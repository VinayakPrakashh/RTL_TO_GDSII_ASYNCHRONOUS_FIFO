* File: pc3b05d.dist.sp
* Created: Sun Jul  4 12:18:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b05d.dist.sp.pex"
.subckt pc3b05d  PAD VSSO VSS VDDO CIN VDD I OEN
* 
M71 N_U29_padr_M71_d N_net_m71_VDDO_res_M71_g U31_U22_source N_VSS_M43_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U31_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M43_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M39 N_PAD_M37_d N_U30_ngate_M39_g N_VSSO_M39_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M37 N_PAD_M37_d N_U29_U42_r1_M37_g N_VSSO_M37_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M40 N_PAD_M41_d N_U30_ngate_M40_g N_VSSO_M40_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M41_d N_U30_ngate_M41_g N_VSSO_M39_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M42_d N_U17_ngate2_M33_g N_VSSO_M33_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M42_d N_U30_ngate_M42_g N_VSSO_M40_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M34 N_PAD_M35_d N_U17_ngate2_M34_g N_VSSO_M34_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M35_d N_U17_ngate2_M35_g N_VSSO_M33_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M31 N_PAD_M36_d N_U29_ngate3_M31_g N_VSSO_M31_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U17_ngate2_M36_g N_VSSO_M34_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M32_d N_U29_U42_r1_M38_g N_VSSO_M38_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M32 N_PAD_M32_d N_U29_ngate3_M32_g N_VSSO_M31_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M44 N_U30_pgate_M44_d N_net_m44_VSSO_res_M44_g N_U29_U72_pgate_M44_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M44@2 N_U30_pgate_M44_d N_net_m44_VSSO_res_M44@2_g N_U29_U72_pgate_M44@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@3 N_U30_pgate_M44@3_d N_net_m44_VSSO_res_M44@3_g N_U29_U72_pgate_M44@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@4 N_U30_pgate_M44@3_d N_net_m44_VSSO_res_M44@4_g N_U29_U72_pgate_M44@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@5 N_U30_pgate_M44@5_d N_net_m44_VSSO_res_M44@5_g N_U29_U72_pgate_M44@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U29_U42_r1_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR45 N_noxref_2_R45_pos N_PAD_R45_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR46 N_noxref_2_R46_pos N_U29_padr_R46_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M59 N_VDDO_M59_d N_U29_U71_UN_P_TOP_M59_g N_PAD_M59_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M60 N_VDDO_M51_d N_U29_U71_UN_P_TOP_M60_g N_PAD_M59_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M49 N_VDDO_M58_d N_U29_U72_pgate_M49_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M50_d N_U29_U72_pgate_M50_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M51 N_VDDO_M51_d N_U29_U72_pgate_M51_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U29_U72_pgate_M52_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U29_U72_pgate_M53_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U29_U72_pgate_M54_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_VDDO_M54_d N_U29_U72_pgate_M55_g N_PAD_M55_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M56 N_VDDO_M56_d N_U29_U72_pgate_M56_g N_PAD_M55_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M57 N_VDDO_M56_d N_U29_U72_pgate_M57_g N_PAD_M57_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M58 N_VDDO_M58_d N_U29_U72_pgate_M58_g N_PAD_M57_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_U30_pgate_M43_d N_net_m43_VDDO_res_M43_g N_U29_U72_pgate_M43_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M43@2 N_U30_pgate_M43_d N_net_m43_VDDO_res_M43@2_g N_U29_U72_pgate_M43@2_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M43@3 N_U30_pgate_M43@3_d N_net_m43_VDDO_res_M43@3_g N_U29_U72_pgate_M43@2_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U29_U71_UN_P_TOP_M62_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M43_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M48 N_U29_ngate3_M48_d N_U17_ngatex_M48_g N_VSSO_M48_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M43_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M43_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M28 N_U30_U12_oenb_M28_d N_U30_U15_OUTSHIFT_M28_g N_VSSO_M28_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M9 N_U30_ngate_M9_d N_U30_ISHF_M9_g N_VSSO_M9_s N_VSS_M43_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M9@2 N_U30_ngate_M9_d N_U30_ISHF_M9@2_g N_VSSO_M9@2_s N_VSS_M43_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M27 N_U30_ngate_M27_d N_U30_U15_OUTSHIFT_M27_g N_VSSO_M9@2_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M10 N_U30_pgate_M10_d N_U30_U12_oenb_M10_g N_U30_ngate_M10_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M10@2 N_U30_pgate_M10@2_d N_U30_U12_oenb_M10@2_g N_U30_ngate_M10_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M10@3 N_U30_pgate_M10@2_d N_U30_U12_oenb_M10@3_g N_U30_ngate_M10@3_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M21 N_U30_U15_MPLL1_dr_M21_d N_OEN_M21_g N_VSSO_M21_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M23 N_VDDO_M23_d N_U30_U15_MN1_drai_M23_g N_U30_U15_MPLL1_dr_M23_s N_VSS_M43_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M21@2 N_U30_U15_MPLL1_dr_M21@2_d N_OEN_M21@2_g N_VSSO_M21_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22 N_U30_U15_OUTSHIFT_M22_d N_U30_U15_MN1_drai_M22_g N_VSSO_M22_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22@2 N_U30_U15_OUTSHIFT_M22@2_d N_U30_U15_MN1_drai_M22@2_g N_VSSO_M22_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M15 N_VDDO_M15_d N_U30_U14_MN1_drai_M15_g N_U30_U14_MPLL1_dr_M15_s N_VSS_M43_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U30_U14_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U30_U14_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U30_ISHF_M14_d N_U30_U14_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U30_ISHF_M14@2_d N_U30_U14_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U30_U14_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M43_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M24 N_U30_U15_MN1_drai_M24_d N_OEN_M24_g N_VSS_M16_s N_VSS_M43_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U29_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M63_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M63_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M47 N_U29_ngate3_M47_d N_U17_ngatex_M47_g N_U17_ngate2_M47_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M29 N_U30_U12_oenb_M29_d N_U30_U15_OUTSHIFT_M29_g N_VDDO_M29_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M29@2 N_U30_U12_oenb_M29@2_d N_U30_U15_OUTSHIFT_M29@2_g N_VDDO_M29_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M7 N_U30_pgate_M7_d N_U30_ISHF_M7_g N_VDDO_M7_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M7@2 N_U30_pgate_M7_d N_U30_ISHF_M7@2_g N_VDDO_M7@2_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M7@3 N_U30_pgate_M7@3_d N_U30_ISHF_M7@3_g N_VDDO_M7@2_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M30 N_U30_pgate_M7@3_d N_U30_U12_oenb_M30_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M30@2 N_U30_pgate_M30@2_d N_U30_U12_oenb_M30@2_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8 N_U30_ngate_M8_d N_U30_U15_OUTSHIFT_M8_g N_U30_pgate_M8_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8@2 N_U30_ngate_M8_d N_U30_U15_OUTSHIFT_M8@2_g N_U30_pgate_M8@2_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_U30_ngate_M8@3_d N_U30_U15_OUTSHIFT_M8@3_g N_U30_pgate_M8@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M19 N_U30_U15_MPLL1_dr_M19_d N_U30_U15_OUTSHIFT_M19_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M20 N_U30_U15_OUTSHIFT_M20_d N_U30_U15_MPLL1_dr_M20_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U30_U14_MPLL1_dr_M11_d N_U30_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U30_ISHF_M12_d N_U30_U14_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M17_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M17 N_U30_U14_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U30_U14_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25 N_U30_U15_MN1_drai_M25_d N_OEN_M25_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25@2 N_U30_U15_MN1_drai_M25_d N_OEN_M25@2_g N_VDD_M25@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D18 N_VSS_M43_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
D26 N_VSS_M43_b N_OEN_D26_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM43 N_VDDO_RM43_pos N_net_m43_VDDO_res_RM43_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM44 N_net_m44_VSSO_res_RM44_pos N_VSSO_RM44_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b05d.dist.sp.PC3B05D.pxi"
*
.ends
*
*
