* File: pt3o01.dist.sp
* Created: Sun Jul  4 13:03:17 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3o01.dist.sp.pex"
.subckt pt3o01  VSS VDDO VSSO I PAD VDD
* 
M29 N_ngate_M29_d N_U28_ISHF_M29_g N_VSSO_M29_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M29@2 N_ngate_M29_d N_U28_ISHF_M29@2_g N_VSSO_M29@2_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M30 N_pgate_M30_d N_net_m30_VDDO_res_M30_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M30@2 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@2_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M30@3 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@3_g N_ngate_M30@3_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_VDDO_M37_d N_U28_U16_MN1_drai_M37_g N_U28_U16_MPLL1_dr_M37_s N_VSS_M29_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M35 N_U28_U16_MPLL1_dr_M35_d N_I_M35_g N_VSSO_M35_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M35@2 N_U28_U16_MPLL1_dr_M35@2_d N_I_M35@2_g N_VSSO_M35_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36 N_U28_ISHF_M36_d N_U28_U16_MN1_drai_M36_g N_VSSO_M36_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36@2 N_U28_ISHF_M36@2_d N_U28_U16_MN1_drai_M36@2_g N_VSSO_M36_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_PAD_M11_d N_U29_U74$9_gate_M5_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M12_d N_U29_U74$9_gate_M6_g N_VSSO_M6_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M13_d N_U29_U74$9_gate_M7_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U29_U74$9_gate_M8_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M3_d N_U29_U74$9_gate_M9_g N_VSSO_M9_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M4_d N_U29_U74$9_gate_M10_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_U28_U16_MN1_drai_M38_d N_I_M38_g N_VSS_M38_s N_VSS_M29_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M31 N_pgate_M31_d N_U28_ISHF_M31_g N_VDDO_M31_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M31@2 N_pgate_M31@2_d N_U28_ISHF_M31@2_g N_VDDO_M31_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M32 N_ngate_M32_d N_net_m32_VSSO_res_M32_g N_pgate_M32_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_ngate_M32_d N_net_m32_VSSO_res_M32@2_g N_pgate_M32@2_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M32@3 N_ngate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_pgate_M32@2_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33 N_U28_U16_MPLL1_dr_M33_d N_U28_ISHF_M33_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M34 N_U28_ISHF_M34_d N_U28_U16_MPLL1_dr_M34_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M39 N_U28_U16_MN1_drai_M39_d N_I_M39_g N_VDD_M39_s N_VDD_M39_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M39@2 N_U28_U16_MN1_drai_M39_d N_I_M39@2_g N_VDD_M39@2_s N_VDD_M39_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D40 N_VSS_M29_b N_I_D40_neg DN18  AREA=2.5e-13 PJ=2e-06
XR27 N_VSSO_R27_pos N_U29_U74$9_gate_R27_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR28 N_U29_U37_r2_R28_pos N_VDDO_R28_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M11 N_PAD_M11_d N_U29_U74$9_gate_M11_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_U74$9_gate_M12_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U74$9_gate_M13_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U29_U74$9_gate_M14_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M3 N_PAD_M3_d N_ngate_M3_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_ngate_M4_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR1 U29_U69_padr N_noxref_11_R1_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR2 N_noxref_11_R2_pos N_PAD_R2_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XRM30 N_net_m30_VDDO_res_RM30_pos N_VDDO_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M17 N_VDDO_M17_d N_U29_U37_r2_M17_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M18 N_VDDO_M19_d N_U29_U37_r2_M18_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M15 N_VDDO_M26_d N_pgate_M15_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M16 N_VDDO_M16_d N_pgate_M16_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M19 N_VDDO_M19_d N_U29_U37_r2_M19_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U29_U37_r2_M20_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U29_U37_r2_M21_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U29_U37_r2_M22_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U29_U37_r2_M23_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U29_U37_r2_M24_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M24_d N_U29_U37_r2_M25_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U37_r2_M26_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U29_U69_padr 0 17.4974f
*
.include "pt3o01.dist.sp.PT3O01.pxi"
*
.ends
*
*
