* File: pvda.dist.sp
* Created: Sun Jul  4 13:18:02 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pvda.dist.sp.pex"
.subckt pvda  VDDO VSSO VSS VDD
* 
M4 N_VDDO_M10_d N_U30_U29_c2_M4_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDO_M11_d N_U30_U29_c2_M5_g N_VSSO_M5_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDO_M12_d N_U30_U29_c2_M6_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_VDDO_M13_d N_U30_U29_c2_M7_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_VDDO_M14_d N_U30_U29_c2_M8_g N_VSSO_M8_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_VDDO_M15_d N_U30_U29_c2_M9_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDO_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U19_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U30_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_VSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_VDDO_M10_d N_U30_U29_c2_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDO_M11_d N_U30_U29_c2_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDO_M12_d N_U30_U29_c2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDO_M13_d N_U30_U29_c2_M13_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDO_M14_d N_U30_U29_c2_M14_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDO_M15_d N_U30_U29_c2_M15_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
D31@2 N_VSSO_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSSO_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSSO_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSSO_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSSO_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSSO_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSSO_D31@8_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSSO_D31@9_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSSO_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@2 N_VSS_D30@2_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSS_D30@3_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSS_D30@4_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSS_D30@5_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSS_D30@6_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSS_D30@7_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSS_D30@8_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSS_D30@9_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSS_D30_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC3_5 N_VDDO_C3_5_pos N_U30_U29_c2_C3_5_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSSO_M16_d N_U19_U22$11_gate_M16_g N_VDDO_M16_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSSO_M16_d N_U19_U22$11_gate_M17_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSSO_M18_d N_U19_U22$11_gate_M18_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSSO_M18_d N_U19_U22$11_gate_M19_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSSO_M20_d N_U19_U22$11_gate_M20_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSSO_M20_d N_U19_U22$11_gate_M21_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSSO_M22_d N_U19_U22$11_gate_M22_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSSO_M22_d N_U19_U22$11_gate_M23_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSSO_M24_d N_U19_U22$11_gate_M24_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSSO_M24_d N_U19_U22$11_gate_M25_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSSO_M26_d N_U19_U22$11_gate_M26_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSSO_M26_d N_U19_U22$11_gate_M27_g N_VDDO_M27_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pvda.dist.sp.PVDA.pxi"
*
.ends
*
*
