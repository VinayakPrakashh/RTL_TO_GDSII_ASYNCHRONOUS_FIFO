* File: pc3d01d.dist.sp
* Created: Sun Jul  4 12:26:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d01d.dist.sp.pex"
.subckt pc3d01d  VSSO VSS VDDO CIN PAD VDD
* 
M1 N_U14_padr_M1_d N_net_m1_VDDO_res_M1_g U15_U22_source N_VSS_M12_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M2 U15_U22_source N_net_m2_VDDO_res_M2_g N_VSSO_M2_s N_VSS_M12_b NHV L=5.5e-06
+ W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M16 N_PAD_M22_d N_U14_MN4$11_gate_M16_g N_VSSO_M16_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M23_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M18 N_PAD_M24_d N_U14_MN4$11_gate_M18_g N_VSSO_M18_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M25_d N_U14_MN4$11_gate_M19_g N_VSSO_M16_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U14_MN4$11_gate_M20_g N_VSSO_M20_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M21 N_PAD_M27_d N_U14_MN4$11_gate_M21_g N_VSSO_M18_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR28 N_U14_MN4$11_gate_R28_pos N_VSSO_R28_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VDDO_res_RM1_pos N_VDDO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_VDDO_RM1_neg N_net_m2_VDDO_res_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
M22 N_PAD_M22_d N_U14_MN4$11_gate_M22_g N_VSSO_M22_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M23_d N_U14_MN4$11_gate_M23_g N_VSSO_M22_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U14_MN4$11_gate_M24_g N_VSSO_M24_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U14_MN4$11_gate_M25_g N_VSSO_M24_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U14_MN4$11_gate_M26_g N_VSSO_M26_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M27 N_PAD_M27_d N_U14_MN4$11_gate_M27_g N_VSSO_M26_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M30 N_VDDO_M33_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M40_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M33 N_VDDO_M33_d N_U14_pgate_tol_M33_g N_PAD_M33_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U14_pgate_tol_M34_g N_PAD_M33_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_VDDO_M34_d N_U14_pgate_tol_M35_g N_PAD_M35_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U14_pgate_tol_M36_g N_PAD_M35_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_VDDO_M36_d N_U14_pgate_tol_M37_g N_PAD_M37_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_VDDO_M38_d N_U14_pgate_tol_M38_g N_PAD_M37_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M39 N_VDDO_M38_d N_U14_pgate_tol_M39_g N_PAD_M39_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M40 N_VDDO_M40_d N_U14_pgate_tol_M40_g N_PAD_M39_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR14 N_X28/noxref_9_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR15 N_X28/noxref_9_R15_pos N_U14_padr_R15_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M12 N_U14_pgate_tol_M12_s N_net_m12_VDDO_res_M12_g N_U14_pgate_tol_M12_s
+ N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M12@2 N_U14_pgate_tol_M12@2_s N_net_m12_VDDO_res_M12@2_g
+ N_U14_pgate_tol_M12@2_s N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M12@3 N_U14_pgate_tol_M12@3_s N_net_m12_VDDO_res_M12@3_g
+ N_U14_pgate_tol_M12@3_s N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M10 N_VDDO_M10_d N_net_m10_VDDO_res_M10_g N_U14_pgate_tol_M10_s N_VSS_M12_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M8 N_U14_padr_M8_d N_net_m8_VSSO_res_M8_g N_VSSO_M8_s N_VSS_M12_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_U14_padr_M8@2_d N_net_m8_VSSO_res_M8@2_g N_VSSO_M8_s N_VSS_M12_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7 N_U9_MPI1_drain_M7_d N_U14_padr_M7_g N_VSSO_M7_s N_VSS_M12_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M9 N_CIN_M9_d N_U9_MPI1_drain_M9_g N_VSS_M9_s N_VSS_M12_b NHV L=3.6e-07 W=6e-06
+ AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M13 N_U14_pgate_tol_M13_s N_net_m13_VSSO_res_M13_g N_U14_pgate_tol_M13_s
+ N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M13@2 N_U14_pgate_tol_M13@2_s N_net_m13_VSSO_res_M13@2_g
+ N_U14_pgate_tol_M13@2_s N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M13@3 N_U14_pgate_tol_M13@3_s N_net_m13_VSSO_res_M13@3_g
+ N_U14_pgate_tol_M13@3_s N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M11 N_U14_pgate_tol_M11_d N_net_m11_VSSO_res_M11_g N_VDDO_M11_s N_VDDO_M13_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M5 N_U14_padr_M5_d N_net_m5_VDDO_res_M5_g N_VDDO_M5_s N_VDDO_M13_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 U9_MPI2_drain N_U14_padr_M3_g N_VDDO_M3_s N_VDDO_M13_b PHV L=3.6e-07 W=2e-05
+ AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M4 N_U9_MPI1_drain_M4_d N_U14_padr_M4_g U9_MPI2_drain N_VDDO_M13_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M6 N_CIN_M6_d N_U9_MPI1_drain_M6_g N_VDD_M6_s N_VDD_M6_b PHV L=3.6e-07 W=8e-06
+ AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M6@2 N_CIN_M6@2_d N_U9_MPI1_drain_M6@2_g N_VDD_M6_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M6@3 N_CIN_M6@2_d N_U9_MPI1_drain_M6@3_g N_VDD_M6@3_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M6@4 N_CIN_M6@4_d N_U9_MPI1_drain_M6@4_g N_VDD_M6@3_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM5 N_net_m5_VDDO_res_RM5_pos N_VDDO_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM13 N_VSSO_RM13_pos N_net_m13_VSSO_res_RM13_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM12 N_VDDO_RM12_pos N_net_m12_VDDO_res_RM12_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM10 N_VDDO_RM10_pos N_net_m10_VDDO_res_RM10_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM11 N_net_m11_VSSO_res_RM11_pos N_VSSO_RM11_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM8 N_VSSO_RM8_pos N_net_m8_VSSO_res_RM8_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U9_MPI2_drain 0 0.0173376f
*
.include "pc3d01d.dist.sp.PC3D01D.pxi"
*
.ends
*
*
