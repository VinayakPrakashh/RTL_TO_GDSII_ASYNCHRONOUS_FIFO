* File: apv0a.dist.sp
* Created: Sun Jul  4 12:04:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apv0a.dist.sp.pex"
.subckt apv0a  AVSSO AVDDO AVSS VSS AVDD
* 
M4 N_AVDDO_M10_d N_U31_U29_c2_M4_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_AVDDO_M11_d N_U31_U29_c2_M5_g N_AVSSO_M5_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_AVDDO_M12_d N_U31_U29_c2_M6_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_AVDDO_M13_d N_U31_U29_c2_M7_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_AVDDO_M14_d N_U31_U29_c2_M8_g N_AVSSO_M8_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_AVDDO_M15_d N_U31_U29_c2_M9_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR16 N_AVDDO_R16_pos N_noxref_3_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR17 N_noxref_3_R17_pos N_U19_U31_r2_R17_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_U31_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_AVSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_AVDDO_M10_d N_U31_U29_c2_M10_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_AVDDO_M11_d N_U31_U29_c2_M11_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_AVDDO_M12_d N_U31_U29_c2_M12_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_AVDDO_M13_d N_U31_U29_c2_M13_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_AVDDO_M14_d N_U31_U29_c2_M14_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_AVDDO_M15_d N_U31_U29_c2_M15_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M18 N_AVSSO_M18_d N_U19_U31_r2_M18_g N_AVDDO_M18_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M19 N_AVSSO_M18_d N_U19_U31_r2_M19_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_AVSSO_M20_d N_U19_U31_r2_M20_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_AVSSO_M20_d N_U19_U31_r2_M21_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_AVSSO_M22_d N_U19_U31_r2_M22_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_AVSSO_M22_d N_U19_U31_r2_M23_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_AVSSO_M24_d N_U19_U31_r2_M24_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_AVSSO_M24_d N_U19_U31_r2_M25_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_AVSSO_M26_d N_U19_U31_r2_M26_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_AVSSO_M26_d N_U19_U31_r2_M27_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M28 N_AVSSO_M28_d N_U19_U31_r2_M28_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M29 N_AVSSO_M28_d N_U19_U31_r2_M29_g N_AVDDO_M29_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
D30@2 N_AVSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_AVSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_AVSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_AVSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_AVSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_AVSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_AVSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_AVSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_AVSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC6_7 N_AVDDO_C6_7_pos N_U31_U29_c2_C6_7_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "apv0a.dist.sp.APV0A.pxi"
*
.ends
*
*
