* File: pc3c01.dist.sp
* Created: Sun Jul  4 12:21:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c01.dist.sp.pex"
.subckt pc3c01  VDD VSS CCLK CP VDDO VSSO
* 
M10 N_NODE_M10_d N_CCLK_M10_g N_VDD_M10_s N_VDD_M10_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M12 N_NODE_M10_d N_CCLK_M12_g N_VDD_M12_s N_VDD_M10_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M4 N_CP_M4_d N_NODE_M4_g N_VDD_M4_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M5 N_CP_M4_d N_NODE_M5_g N_VDD_M5_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M8 N_CP_M8_d N_NODE_M8_g N_VDD_M5_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M9 N_CP_M8_d N_NODE_M9_g N_VDD_M9_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D1 N_VSS_M11_b N_CCLK_D1_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M11 N_NODE_M11_d N_CCLK_M11_g N_VSS_M11_s N_VSS_M11_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M13 N_NODE_M11_d N_CCLK_M13_g N_VSS_M13_s N_VSS_M11_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M2 N_CP_M2_d N_NODE_M2_g N_VSS_M2_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M3 N_CP_M2_d N_NODE_M3_g N_VSS_M3_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_CP_M6_d N_NODE_M6_g N_VSS_M3_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M7 N_CP_M6_d N_NODE_M7_g N_VSS_M7_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
*
.include "pc3c01.dist.sp.PC3C01.pxi"
*
.ends
*
*
