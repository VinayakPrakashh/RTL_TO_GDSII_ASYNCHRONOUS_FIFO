* File: pc3d21.dist.sp
* Created: Sun Jul  4 12:31:01 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d21.dist.sp.pex"
.subckt pc3d21  VSS VSSO CIN PAD VDDO VDD
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X24/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X24/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U14_padr_M34_d N_net_m34_VSSO_res_M34_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M34@2 N_U14_padr_M34@2_d N_net_m34_VSSO_res_M34@2_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M32 N_U9_U34_drain_M32_d N_U14_padr_M32_g N_VSSO_M32_s N_VSS_M3_b NHV L=3.6e-07
+ W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M33 N_U9_U36_drain_M33_d N_U14_padr_M33_g N_U9_U34_drain_M32_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M35 N_VDDO_M35_d N_U9_U36_drain_M35_g N_U9_U34_drain_M35_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M36 N_CIN_M36_d N_U9_U36_drain_M36_g N_VSS_M36_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M39 N_U14_padr_M39_d N_net_m39_VDDO_res_M39_g N_VDDO_M39_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M39@2 N_U14_padr_M39_d N_net_m39_VDDO_res_M39@2_g N_VDDO_M39@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38 N_U9_U30_source_M38_d N_U14_padr_M38_g N_VDDO_M38_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M37 N_U9_U36_drain_M37_d N_U14_padr_M37_g N_U9_U30_source_M38_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M40 N_VSSO_M40_d N_U9_U36_drain_M40_g N_U9_U30_source_M40_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M41 N_CIN_M41_d N_U9_U36_drain_M41_g N_VDD_M41_s N_VDD_M41_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M41@2 N_CIN_M41@2_d N_U9_U36_drain_M41@2_g N_VDD_M41_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@3 N_CIN_M41@2_d N_U9_U36_drain_M41@3_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@4 N_CIN_M41@4_d N_U9_U36_drain_M41@4_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM39 N_net_m39_VDDO_res_RM39_pos N_VDDO_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM34 N_VSSO_RM34_pos N_net_m34_VSSO_res_RM34_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d21.dist.sp.PC3D21.pxi"
*
.ends
*
*
