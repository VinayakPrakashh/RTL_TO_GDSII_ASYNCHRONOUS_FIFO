* File: pc3t02.dist.sp
* Created: Sun Jul  4 12:43:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t02.dist.sp.pex"
.subckt pc3t02  PAD VSS VSSO VDDO VDD I OEN
* 
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M65 N_U27_padr_M65_d N_net_m65_VSSO_res_M65_g N_VSSO_M65_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M65@2 N_U27_padr_M65@2_d N_net_m65_VSSO_res_M65@2_g N_VSSO_M65_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U28_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U28_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U28_MPI1_drain_M63_d N_U27_padr_M63_g U28_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM65 N_VSSO_RM65_pos N_net_m65_VSSO_res_RM65_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.361103f
c_2 U28_MPI2_drain 0 0.0169448f
*
.include "pc3t02.dist.sp.PC3T02.pxi"
*
.ends
*
*
