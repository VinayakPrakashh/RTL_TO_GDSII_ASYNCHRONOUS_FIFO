/run/media/user1/c2s/S5_training_batch2/VINAYAK/05_Floorplanning/tsl180l4.lef