* File: pc3c04.dist.sp
* Created: Sun Jul  4 12:24:16 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c04.dist.sp.pex"
.subckt pc3c04  CCLK VDD CP VSS VDDO VSSO
* 
M1 N_CP_M33_d N_NODE_M1_g N_VSS_M1_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M2 N_CP_M34_d N_NODE_M2_g N_VSS_M2_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M5 N_CP_M37_d N_NODE_M5_g N_VSS_M2_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_CP_M38_d N_NODE_M6_g N_VSS_M6_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M9 N_CP_M41_d N_NODE_M9_g N_VSS_M6_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M10 N_CP_M42_d N_NODE_M10_g N_VSS_M10_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M13 N_CP_M45_d N_NODE_M13_g N_VSS_M10_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_CP_M46_d N_NODE_M14_g N_VSS_M14_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M17 N_CP_M49_d N_NODE_M17_g N_VSS_M14_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M18 N_CP_M50_d N_NODE_M18_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M21 N_CP_M53_d N_NODE_M21_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M54_d N_NODE_M22_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M25 N_CP_M57_d N_NODE_M25_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M26 N_CP_M58_d N_NODE_M26_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M29 N_CP_M61_d N_NODE_M29_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M30 N_CP_M62_d N_NODE_M30_g N_VSS_M30_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M65 N_NODE_M65_d N_CCLK_M65_g N_VDD_M65_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M67 N_NODE_M65_d N_CCLK_M67_g N_VDD_M67_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M69 N_NODE_M69_d N_CCLK_M69_g N_VDD_M69_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M71 N_NODE_M69_d N_CCLK_M71_g N_VDD_M71_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M73 N_NODE_M73_d N_CCLK_M73_g N_VDD_M73_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M75 N_NODE_M73_d N_CCLK_M75_g N_VDD_M75_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M77 N_NODE_M77_d N_CCLK_M77_g N_VDD_M77_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M79 N_NODE_M77_d N_CCLK_M79_g N_VDD_M79_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M81 N_NODE_M81_d N_CCLK_M81_g N_VDD_M81_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M83 N_NODE_M81_d N_CCLK_M83_g N_VDD_M83_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M85 N_NODE_M85_d N_CCLK_M85_g N_VDD_M85_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M87 N_NODE_M85_d N_CCLK_M87_g N_VDD_M87_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M89 N_NODE_M89_d N_CCLK_M89_g N_VDD_M89_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M91 N_NODE_M89_d N_CCLK_M91_g N_VDD_M91_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M93 N_NODE_M93_d N_CCLK_M93_g N_VDD_M93_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M95 N_NODE_M93_d N_CCLK_M95_g N_VDD_M95_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_CP_M3_d N_NODE_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M4 N_CP_M3_d N_NODE_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M7 N_CP_M7_d N_NODE_M7_g N_VDD_M4_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M8 N_CP_M7_d N_NODE_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M11 N_CP_M11_d N_NODE_M11_g N_VDD_M8_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M12 N_CP_M11_d N_NODE_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M15 N_CP_M15_d N_NODE_M15_g N_VDD_M12_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M16 N_CP_M15_d N_NODE_M16_g N_VDD_M16_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M16_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M27 N_CP_M27_d N_NODE_M27_g N_VDD_M24_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M28 N_CP_M27_d N_NODE_M28_g N_VDD_M28_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M31 N_CP_M31_d N_NODE_M31_g N_VDD_M28_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M32 N_CP_M31_d N_NODE_M32_g N_VDD_M32_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M35 N_CP_M35_d N_NODE_M35_g N_VDD_M32_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M36 N_CP_M35_d N_NODE_M36_g N_VDD_M36_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M39 N_CP_M39_d N_NODE_M39_g N_VDD_M36_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M40 N_CP_M39_d N_NODE_M40_g N_VDD_M40_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M43 N_CP_M43_d N_NODE_M43_g N_VDD_M40_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M44 N_CP_M43_d N_NODE_M44_g N_VDD_M44_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M47 N_CP_M47_d N_NODE_M47_g N_VDD_M44_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M48 N_CP_M47_d N_NODE_M48_g N_VDD_M48_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M51 N_CP_M51_d N_NODE_M51_g N_VDD_M48_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M52 N_CP_M51_d N_NODE_M52_g N_VDD_M52_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M55 N_CP_M55_d N_NODE_M55_g N_VDD_M52_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M56 N_CP_M55_d N_NODE_M56_g N_VDD_M56_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M59 N_CP_M59_d N_NODE_M59_g N_VDD_M56_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M60 N_CP_M59_d N_NODE_M60_g N_VDD_M60_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M63 N_CP_M63_d N_NODE_M63_g N_VDD_M60_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M64 N_CP_M63_d N_NODE_M64_g N_VDD_M64_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D97 N_VSS_M66_b N_CCLK_D97_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M66 N_NODE_M66_d N_CCLK_M66_g N_VSS_M66_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M68 N_NODE_M66_d N_CCLK_M68_g N_VSS_M68_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M33 N_CP_M33_d N_NODE_M33_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M34 N_CP_M34_d N_NODE_M34_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M70 N_NODE_M70_d N_CCLK_M70_g N_VSS_M70_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M72 N_NODE_M70_d N_CCLK_M72_g N_VSS_M72_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_CP_M37_d N_NODE_M37_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M38 N_CP_M38_d N_NODE_M38_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M74 N_NODE_M74_d N_CCLK_M74_g N_VSS_M74_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M76 N_NODE_M74_d N_CCLK_M76_g N_VSS_M76_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41 N_CP_M41_d N_NODE_M41_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M42 N_CP_M42_d N_NODE_M42_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M78 N_NODE_M78_d N_CCLK_M78_g N_VSS_M78_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M80 N_NODE_M78_d N_CCLK_M80_g N_VSS_M80_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_CP_M45_d N_NODE_M45_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M46 N_CP_M46_d N_NODE_M46_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M82 N_NODE_M82_d N_CCLK_M82_g N_VSS_M82_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M84 N_NODE_M82_d N_CCLK_M84_g N_VSS_M84_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M49 N_CP_M49_d N_NODE_M49_g N_VSS_M49_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M50 N_CP_M50_d N_NODE_M50_g N_VSS_M49_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M86 N_NODE_M86_d N_CCLK_M86_g N_VSS_M86_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M88 N_NODE_M86_d N_CCLK_M88_g N_VSS_M88_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M53 N_CP_M53_d N_NODE_M53_g N_VSS_M53_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M54 N_CP_M54_d N_NODE_M54_g N_VSS_M53_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M90 N_NODE_M90_d N_CCLK_M90_g N_VSS_M90_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M92 N_NODE_M90_d N_CCLK_M92_g N_VSS_M92_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M57 N_CP_M57_d N_NODE_M57_g N_VSS_M57_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M58 N_CP_M58_d N_NODE_M58_g N_VSS_M57_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M94 N_NODE_M94_d N_CCLK_M94_g N_VSS_M94_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M96 N_NODE_M94_d N_CCLK_M96_g N_VSS_M96_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M61 N_CP_M61_d N_NODE_M61_g N_VSS_M61_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M62 N_CP_M62_d N_NODE_M62_g N_VSS_M61_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c04.dist.sp.PC3C04.pxi"
*
.ends
*
*
