* File: pc3d00.dist.sp
* Created: Sun Jul  4 12:24:11 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d00.dist.sp.pex"
.subckt pc3d00  PADR PAD VSS VDDO VSSO VDD
* 
M19 N_PAD_M25_d N_U18_U74$11_gate_M19_g N_VSSO_M19_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U18_U74$11_gate_M20_g N_VSSO_M20_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M21 N_PAD_M27_d N_U18_U74$11_gate_M21_g N_VSSO_M21_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M22 N_PAD_M28_d N_U18_U74$11_gate_M22_g N_VSSO_M19_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M29_d N_U18_U74$11_gate_M23_g N_VSSO_M23_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M24 N_PAD_M30_d N_U18_U74$11_gate_M24_g N_VSSO_M21_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
D32@2 N_VSS_D32@2_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@3 N_VSS_D32@3_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@4 N_VSS_D32@4_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@5 N_VSS_D32@5_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@6 N_VSS_D32@6_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@7 N_VSS_D32@7_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32 N_VSS_D32_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSSO_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSSO_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSSO_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSSO_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSSO_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSSO_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSSO_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XR15 N_VSS_R15_pos N_U18_U82_gate_R15_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR16 N_U18_U74$11_gate_R16_pos N_VSSO_R16_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR17 N_U18_U79$3_gate_R17_pos N_VDDO_R17_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M25 N_PAD_M25_d N_U18_U74$11_gate_M25_g N_VSSO_M25_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U18_U74$11_gate_M26_g N_VSSO_M25_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M27 N_PAD_M27_d N_U18_U74$11_gate_M27_g N_VSSO_M27_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M28 N_PAD_M28_d N_U18_U74$11_gate_M28_g N_VSSO_M27_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M29 N_PAD_M29_d N_U18_U74$11_gate_M29_g N_VSSO_M29_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M30 N_PAD_M30_d N_U18_U74$11_gate_M30_g N_VSSO_M29_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR13 N_PADR_R13_pos N_noxref_2_R13_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR14 N_noxref_2_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M1 N_VDDO_M1_d N_U18_U79$3_gate_M1_g N_PAD_M1_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M2 N_VDDO_M5_d N_U18_U79$3_gate_M2_g N_PAD_M1_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_VDDO_M12_d N_U18_U79$3_gate_M3_g N_PAD_M3_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M4 N_VDDO_M4_d N_U18_U79$3_gate_M4_g N_PAD_M3_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M5 N_VDDO_M5_d N_U18_U79$3_gate_M5_g N_PAD_M5_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M6 N_VDDO_M6_d N_U18_U79$3_gate_M6_g N_PAD_M5_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M7 N_VDDO_M6_d N_U18_U79$3_gate_M7_g N_PAD_M7_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M8 N_VDDO_M8_d N_U18_U79$3_gate_M8_g N_PAD_M7_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M9 N_VDDO_M8_d N_U18_U79$3_gate_M9_g N_PAD_M9_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M10 N_VDDO_M10_d N_U18_U79$3_gate_M10_g N_PAD_M9_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M11 N_VDDO_M10_d N_U18_U79$3_gate_M11_g N_PAD_M11_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M12 N_VDDO_M12_d N_U18_U79$3_gate_M12_g N_PAD_M11_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_PADR_M18_d N_U18_U82_gate_M18_g N_VSS_M18_s N_VSS_M18_b NHV L=4e-07
+ W=3e-05 AD=1.842e-10 AS=4.29e-11 PD=7.228e-05 PS=6.286e-05
*
.include "pc3d00.dist.sp.PC3D00.pxi"
*
.ends
*
*
