* File: apc3d01.dist.sp
* Created: Sun Jul  4 12:03:25 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apc3d01.dist.sp.pex"
.subckt apc3d01  PAD CIN AVSS AVSSO AVDDO AVDD VSS
* 
M7 N_CIN_M7_d N_U9_MPI1_drain_M7_g N_AVSS_M7_s N_AVSS_M7_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M15 N_PAD_M21_d N_U14_U71_r1_M15_g N_AVSSO_M15_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M22_d N_U14_U71_r1_M16_g N_AVSSO_M16_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M17 N_PAD_M23_d N_U14_U71_r1_M17_g N_AVSSO_M17_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M24_d N_U14_U71_r1_M18_g N_AVSSO_M15_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M25_d N_U14_U71_r1_M19_g N_AVSSO_M19_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M20 N_PAD_M26_d N_U14_U71_r1_M20_g N_AVSSO_M17_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR8 N_U14_U71_r1_R8_pos N_AVSSO_R8_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M21 N_PAD_M21_d N_U14_U71_r1_M21_g N_AVSSO_M21_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M22 N_PAD_M22_d N_U14_U71_r1_M22_g N_AVSSO_M21_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M23_d N_U14_U71_r1_M23_g N_AVSSO_M23_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U14_U71_r1_M24_g N_AVSSO_M23_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U14_U71_r1_M25_g N_AVSSO_M25_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U14_U71_r1_M26_g N_AVSSO_M25_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR11 N_PAD_R11_pos N_noxref_2_R11_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR12 N_noxref_2_R12_pos N_U14_padr_R12_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M27 N_AVDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M27_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M28 N_AVDDO_M31_d N_U14_pgate_tol_M28_g N_PAD_M27_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_AVDDO_M38_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_AVDDO_M30_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M31 N_AVDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_AVDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_AVDDO_M32_d N_U14_pgate_tol_M33_g N_PAD_M33_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_AVDDO_M34_d N_U14_pgate_tol_M34_g N_PAD_M33_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_AVDDO_M34_d N_U14_pgate_tol_M35_g N_PAD_M35_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_AVDDO_M36_d N_U14_pgate_tol_M36_g N_PAD_M35_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_AVDDO_M36_d N_U14_pgate_tol_M37_g N_PAD_M37_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_AVDDO_M38_d N_U14_pgate_tol_M38_g N_PAD_M37_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M9 N_U14_pgate_tol_M9_s N_net_m9_AVDDO_res_M9_g N_U14_pgate_tol_M9_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M9@2 N_U14_pgate_tol_M9@2_s N_net_m9_AVDDO_res_M9@2_g N_U14_pgate_tol_M9@2_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M9@3 N_U14_pgate_tol_M9@3_s N_net_m9_AVDDO_res_M9@3_g N_U14_pgate_tol_M9@3_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M13 N_AVDDO_M13_d N_net_m13_AVDDO_res_M13_g N_U14_pgate_tol_M13_s N_AVSSO_M9_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M6 N_U14_padr_M6_d N_net_m6_AVSSO_res_M6_g N_AVSSO_M6_s N_AVSSO_M9_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6@2 N_U14_padr_M6@2_d N_net_m6_AVSSO_res_M6@2_g N_AVSSO_M6_s N_AVSSO_M9_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_U9_MPI1_drain_M5_d N_U14_padr_M5_g N_AVSSO_M5_s N_AVSSO_M9_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M14 N_U14_pgate_tol_M14_d N_net_m14_AVSSO_res_M14_g N_AVDDO_M14_s N_AVDDO_M14_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 N_U14_padr_M3_d N_net_m3_AVDDO_res_M3_g N_AVDDO_M3_s N_AVDDO_M14_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M1 U9_MPI2_drain N_U14_padr_M1_g N_AVDDO_M1_s N_AVDDO_M14_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M2 N_U9_MPI1_drain_M2_d N_U14_padr_M2_g U9_MPI2_drain N_AVDDO_M14_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M10 N_U14_pgate_tol_M10_s N_net_m10_AVSSO_res_M10_g N_U14_pgate_tol_M10_s
+ N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M10@2 N_U14_pgate_tol_M10@2_s N_net_m10_AVSSO_res_M10@2_g
+ N_U14_pgate_tol_M10@2_s N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M10@3 N_U14_pgate_tol_M10@3_s N_net_m10_AVSSO_res_M10@3_g
+ N_U14_pgate_tol_M10@3_s N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M4 N_CIN_M4_d N_U9_MPI1_drain_M4_g N_AVDD_M4_s N_AVDD_M4_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M4@2 N_CIN_M4@2_d N_U9_MPI1_drain_M4@2_g N_AVDD_M4_s N_AVDD_M4_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M4@3 N_CIN_M4@2_d N_U9_MPI1_drain_M4@3_g N_AVDD_M4@3_s N_AVDD_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M4@4 N_CIN_M4@4_d N_U9_MPI1_drain_M4@4_g N_AVDD_M4@3_s N_AVDD_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
D40@2 N_VSS_D40@2_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@3 N_VSS_D40@3_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@4 N_VSS_D40@4_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@5 N_VSS_D40@5_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@6 N_VSS_D40@6_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@7 N_VSS_D40@7_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40 N_VSS_D40_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@2 N_AVSSO_D39@2_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@3 N_AVSSO_D39@3_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@4 N_AVSSO_D39@4_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@5 N_AVSSO_D39@5_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@6 N_AVSSO_D39@6_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@7 N_AVSSO_D39@7_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39 N_AVSSO_D39_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XRM14 N_AVSSO_RM14_pos N_net_m14_AVSSO_res_RM14_neg RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM3 N_net_m3_AVDDO_res_RM3_pos N_AVDDO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM10 N_AVSSO_RM10_pos N_net_m10_AVSSO_res_RM10_neg RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM9 N_AVDDO_RM9_pos N_net_m9_AVDDO_res_RM9_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM13 N_net_m13_AVDDO_res_RM13_pos N_AVDDO_RM9_pos RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM6 N_net_m6_AVSSO_res_RM6_pos N_AVSSO_RM6_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U9_MPI2_drain 0 0.0183971f
*
.include "apc3d01.dist.sp.APC3D01.pxi"
*
.ends
*
*
