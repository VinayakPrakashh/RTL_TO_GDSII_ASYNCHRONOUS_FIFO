/run/media/user1/c2s/cadence/install/SCLPDK/scl_pdk/stdlib/fs120/lef/tsl18fs120_scl.lef