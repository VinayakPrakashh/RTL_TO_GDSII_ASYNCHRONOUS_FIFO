* File: pt3t01.dist.sp
* Created: Sun Jul  4 13:05:03 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t01.dist.sp.pex"
.subckt pt3t01  PAD VSS VSSO VDDO VDD I OEN
* 
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M59 N_U27_padr_M59_d N_net_m59_VSSO_res_M59_g N_VSSO_M59_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M59@2 N_U27_padr_M59@2_d N_net_m59_VSSO_res_M59@2_g N_VSSO_M59_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60 N_U28_MPI1_drain_M60_d N_U27_padr_M60_g N_VSSO_M60_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 N_U27_padr_M58_d N_net_m58_VDDO_res_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M56 U28_MPI2_drain N_U27_padr_M56_g N_VDDO_M56_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M57 N_U28_MPI1_drain_M57_d N_U27_padr_M57_g U28_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM58 N_net_m58_VDDO_res_RM58_pos N_VDDO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM59 N_VSSO_RM59_pos N_net_m59_VSSO_res_RM59_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U28_MPI2_drain 0 0.0289375f
*
.include "pt3t01.dist.sp.PT3T01.pxi"
*
.ends
*
*
