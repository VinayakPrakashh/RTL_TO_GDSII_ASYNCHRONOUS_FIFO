* File: pt3o03.dist.sp
* Created: Sun Jul  4 13:05:17 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3o03.dist.sp.pex"
.subckt pt3o03  PAD VSS VDDO VSSO I VDD
* 
M13 N_PAD_M15_d N_ngate_M13_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M16_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M9_d N_U30_ngate2_M7_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M10_d N_ngate_M14_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M11_d N_U29_U76_r1_M18_g N_VSSO_M18_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M12_d N_U30_ngate2_M8_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M15 N_PAD_M15_d N_ngate_M15_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_ngate_M16_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M9_d N_U30_ngate2_M9_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U30_ngate2_M10_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U29_ngate3_M11_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_ngate3_M12_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 U29_U69_padr N_noxref_2_R19_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR20 N_noxref_2_R20_pos N_PAD_R20_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M33 N_VDDO_M33_d N_U29_U37_r2_M33_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M25_d N_U29_U37_r2_M34_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_pgate_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_pgate_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_pgate_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_pgate_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_pgate_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_pgate_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_pgate_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_pgate_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M22 N_U29_ngate3_M22_d N_U30_ngatex_M22_g N_VSSO_M22_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U27_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U27_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U27_U13_MN1_drai_M45_g N_U27_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U27_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U27_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U27_ISHF_M44_d N_U27_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U27_ISHF_M44@2_d N_U27_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U27_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M21 N_U29_ngate3_M21_d N_U30_ngatex_M21_g N_U30_ngate2_M21_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U27_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U27_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U27_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U27_U13_MPLL1_dr_M41_d N_U27_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U27_ISHF_M42_d N_U27_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U27_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U27_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.4884f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pt3o03.dist.sp.PT3O03.pxi"
*
.ends
*
*
