* File: pc3c02.dist.sp
* Created: Sun Jul  4 12:22:40 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c02.dist.sp.pex"
.subckt pc3c02  VSS VDD CCLK CP VDDO VSSO
* 
M1 N_NODE_M1_d N_CCLK_M1_g N_VDD_M1_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_NODE_M1_d N_CCLK_M3_g N_VDD_M3_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M5 N_NODE_M5_d N_CCLK_M5_g N_VDD_M5_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M7 N_NODE_M5_d N_CCLK_M7_g N_VDD_M7_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M11 N_CP_M11_d N_NODE_M11_g N_VDD_M11_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M12 N_CP_M11_d N_NODE_M12_g N_VDD_M12_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M15 N_CP_M15_d N_NODE_M15_g N_VDD_M12_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M16 N_CP_M15_d N_NODE_M16_g N_VDD_M16_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M16_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D25 N_VSS_M2_b N_CCLK_D25_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M9 N_CP_M17_d N_NODE_M9_g N_VSS_M9_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M10 N_CP_M18_d N_NODE_M10_g N_VSS_M10_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M13 N_CP_M21_d N_NODE_M13_g N_VSS_M10_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_CP_M22_d N_NODE_M14_g N_VSS_M14_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M2 N_NODE_M2_d N_CCLK_M2_g N_VSS_M2_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4 N_NODE_M2_d N_CCLK_M4_g N_VSS_M4_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M17 N_CP_M17_d N_NODE_M17_g N_VSS_M17_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M18 N_CP_M18_d N_NODE_M18_g N_VSS_M17_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_NODE_M6_d N_CCLK_M6_g N_VSS_M6_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8 N_NODE_M6_d N_CCLK_M8_g N_VSS_M8_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M21 N_CP_M21_d N_NODE_M21_g N_VSS_M21_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M22_d N_NODE_M22_g N_VSS_M21_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c02.dist.sp.PC3C02.pxi"
*
.ends
*
*
