* File: pc3t01.dist.sp
* Created: Sun Jul  4 12:40:31 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t01.dist.sp.pex"
.subckt pc3t01  PAD VSS VSSO VDDO VDD I OEN
* 
M32 N_PAD_M33_d N_U27_U69$9_gate_M32_g N_VSSO_M32_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M33_d N_U27_U69$9_gate_M33_g N_VSSO_M33_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M35_d N_U27_U69$9_gate_M34_g N_VSSO_M34_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M35_d N_U27_U69$9_gate_M35_g N_VSSO_M32_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M37_d N_U27_U69$9_gate_M36_g N_VSSO_M36_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M37 N_PAD_M37_d N_U27_U69$9_gate_M37_g N_VSSO_M34_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M39_d N_U27_U69$9_gate_M38_g N_VSSO_M38_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M39 N_PAD_M39_d N_U27_U69$9_gate_M39_g N_VSSO_M36_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M30 N_PAD_M40_d N_U15_ngate_M30_g N_VSSO_M30_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U27_U69$9_gate_M40_g N_VSSO_M38_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M31_d N_U27_U69$9_gate_M41_g N_VSSO_M41_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M31 N_PAD_M31_d N_U15_ngate_M31_g N_VSSO_M30_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M55 N_U15_pgate_M55_d N_net_m55_VSSO_res_M55_g N_U27_U72_pgate_M55_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M55@2 N_U15_pgate_M55_d N_net_m55_VSSO_res_M55@2_g N_U27_U72_pgate_M55@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@3 N_U15_pgate_M55@3_d N_net_m55_VSSO_res_M55@3_g N_U27_U72_pgate_M55@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@4 N_U15_pgate_M55@3_d N_net_m55_VSSO_res_M55@4_g N_U27_U72_pgate_M55@4_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@5 N_U15_pgate_M55@5_d N_net_m55_VSSO_res_M55@5_g N_U27_U72_pgate_M55@4_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR58 N_U27_U69$9_gate_R58_pos N_VSSO_R58_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR56 N_noxref_2_R56_pos N_PAD_R56_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR57 N_noxref_2_R57_pos N_U27_padr_R57_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M44 N_VDDO_M44_d N_U27_U71_UN_P_TOP_M44_g N_PAD_M44_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M45 N_VDDO_M46_d N_U27_U71_UN_P_TOP_M45_g N_PAD_M44_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M42 N_VDDO_M53_d N_U27_U72_pgate_M42_g N_PAD_M42_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M43_d N_U27_U72_pgate_M43_g N_PAD_M42_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M46 N_VDDO_M46_d N_U27_U71_UN_P_TOP_M46_g N_PAD_M46_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M47 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M47_g N_PAD_M46_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M48 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M48_g N_PAD_M48_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M49 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M49_g N_PAD_M48_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M50_g N_PAD_M50_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M51 N_VDDO_M51_d N_U27_U71_UN_P_TOP_M51_g N_PAD_M50_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M51_d N_U27_U71_UN_P_TOP_M52_g N_PAD_M52_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M53_d N_U27_U71_UN_P_TOP_M53_g N_PAD_M52_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_U15_pgate_M54_d N_net_m54_VDDO_res_M54_g N_U27_U72_pgate_M54_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M54@2 N_U15_pgate_M54_d N_net_m54_VDDO_res_M54@2_g N_U27_U72_pgate_M54@2_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M54@3 N_U15_pgate_M54@3_d N_net_m54_VDDO_res_M54@3_g N_U27_U72_pgate_M54@2_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M59 N_VDDO_M59_d N_net_m59_VDDO_res_M59_g N_U27_U71_UN_P_TOP_M59_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M4 N_U27_padr_M4_d N_net_m4_VSSO_res_M4_g N_VSSO_M4_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M4@2 N_U27_padr_M4@2_d N_net_m4_VSSO_res_M4@2_g N_VSSO_M4_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_U28_MPI1_drain_M5_d N_U27_padr_M5_g N_VSSO_M5_s N_VSS_M54_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M27 N_U15_U12_oenb_M27_d N_U15_U15_OUTSHIFT_M27_g N_VSSO_M27_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M6 N_U15_ngate_M6_d N_U15_ISHF_M6_g N_VSSO_M6_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M6@2 N_U15_ngate_M6_d N_U15_ISHF_M6@2_g N_VSSO_M6@2_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M26 N_U15_ngate_M26_d N_U15_U15_OUTSHIFT_M26_g N_VSSO_M6@2_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M7 N_U15_pgate_M7_d N_U15_U12_oenb_M7_g N_U15_ngate_M7_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7@2 N_U15_pgate_M7@2_d N_U15_U12_oenb_M7@2_g N_U15_ngate_M7_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M7@3 N_U15_pgate_M7@2_d N_U15_U12_oenb_M7@3_g N_U15_ngate_M7@3_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M20 N_U15_U15_MPLL1_dr_M20_d N_OEN_M20_g N_VSSO_M20_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M22 N_VDDO_M22_d N_U15_U15_MN1_drai_M22_g N_U15_U15_MPLL1_dr_M22_s N_VSS_M54_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M20@2 N_U15_U15_MPLL1_dr_M20@2_d N_OEN_M20@2_g N_VSSO_M20_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M21 N_U15_U15_OUTSHIFT_M21_d N_U15_U15_MN1_drai_M21_g N_VSSO_M21_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M21@2 N_U15_U15_OUTSHIFT_M21@2_d N_U15_U15_MN1_drai_M21@2_g N_VSSO_M21_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M14 N_VDDO_M14_d N_U15_U14_MN1_drai_M14_g N_U15_U14_MPLL1_dr_M14_s N_VSS_M54_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M12 N_U15_U14_MPLL1_dr_M12_d N_I_M12_g N_VSSO_M12_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M12@2 N_U15_U14_MPLL1_dr_M12@2_d N_I_M12@2_g N_VSSO_M12_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13 N_U15_ISHF_M13_d N_U15_U14_MN1_drai_M13_g N_VSSO_M13_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U15_ISHF_M13@2_d N_U15_U14_MN1_drai_M13@2_g N_VSSO_M13_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M15 N_U15_U14_MN1_drai_M15_d N_I_M15_g N_VSS_M15_s N_VSS_M54_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M23 N_U15_U15_MN1_drai_M23_d N_OEN_M23_g N_VSS_M15_s N_VSS_M54_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M60 N_U27_U71_UN_P_TOP_M60_d N_net_m60_VSSO_res_M60_g N_VDDO_M60_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 N_U27_padr_M3_d N_net_m3_VDDO_res_M3_g N_VDDO_M3_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M1 U28_MPI2_drain N_U27_padr_M1_g N_VDDO_M1_s N_VDDO_M60_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M2 N_U28_MPI1_drain_M2_d N_U27_padr_M2_g U28_MPI2_drain N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M28 N_U15_U12_oenb_M28_d N_U15_U15_OUTSHIFT_M28_g N_VDDO_M28_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M28@2 N_U15_U12_oenb_M28@2_d N_U15_U15_OUTSHIFT_M28@2_g N_VDDO_M28_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M8 N_U15_pgate_M8_d N_U15_ISHF_M8_g N_VDDO_M8_s N_VDDO_M60_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M8@2 N_U15_pgate_M8@2_d N_U15_ISHF_M8@2_g N_VDDO_M8_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M29 N_U15_pgate_M8@2_d N_U15_U12_oenb_M29_g N_VDDO_M29_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M29@2 N_U15_pgate_M29@2_d N_U15_U12_oenb_M29@2_g N_VDDO_M29_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M9 N_U15_ngate_M9_d N_U15_U15_OUTSHIFT_M9_g N_U15_pgate_M9_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9@2 N_U15_ngate_M9_d N_U15_U15_OUTSHIFT_M9@2_g N_U15_pgate_M9@2_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M9@3 N_U15_ngate_M9@3_d N_U15_U15_OUTSHIFT_M9@3_g N_U15_pgate_M9@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M18 N_U15_U15_MPLL1_dr_M18_d N_U15_U15_OUTSHIFT_M18_g N_VDDO_M18_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M19 N_U15_U15_OUTSHIFT_M19_d N_U15_U15_MPLL1_dr_M19_g N_VDDO_M18_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M10 N_U15_U14_MPLL1_dr_M10_d N_U15_ISHF_M10_g N_VDDO_M10_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U15_ISHF_M11_d N_U15_U14_MPLL1_dr_M11_g N_VDDO_M10_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M16 N_U15_U14_MN1_drai_M16_d N_I_M16_g N_VDD_M16_s N_VDD_M16_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M16@2 N_U15_U14_MN1_drai_M16_d N_I_M16@2_g N_VDD_M16@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M24 N_U15_U15_MN1_drai_M24_d N_OEN_M24_g N_VDD_M16@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M24@2 N_U15_U15_MN1_drai_M24_d N_OEN_M24@2_g N_VDD_M24@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D17 N_VSS_M54_b N_I_D17_neg DN18  AREA=2.5e-13 PJ=2e-06
D25 N_VSS_M54_b N_OEN_D25_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM60 N_VSSO_RM60_pos N_net_m60_VSSO_res_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM3 N_net_m3_VDDO_res_RM3_pos N_VDDO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM54 N_VDDO_RM54_pos N_net_m54_VDDO_res_RM54_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM59 N_VDDO_RM59_pos N_net_m59_VDDO_res_RM59_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM55 N_net_m55_VSSO_res_RM55_pos N_VSSO_RM55_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U28_MPI2_drain 0 0.0289375f
*
.include "pc3t01.dist.sp.PC3T01.pxi"
*
.ends
*
*
