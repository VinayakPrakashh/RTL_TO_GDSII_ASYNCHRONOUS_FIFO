* File: pv0c.dist.sp
* Created: Sun Jul  4 13:13:03 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0c.dist.sp.pex"
.subckt pv0c  VSSC VDD VDDO VSS VSSO
* 
M18 N_VDD_M19_d N_U33_U29_c2_M18_g N_VSSC_M25_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_VDD_M19_d N_U33_U29_c2_M19_g N_VSSC_M19_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_VDD_M21_d N_U33_U29_c2_M20_g N_VSSC_M20_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M21 N_VDD_M21_d N_U33_U29_c2_M21_g N_VSSC_M26_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_VDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U34_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_U33_U29_c2_R16_pos N_noxref_7_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR17 N_noxref_7_R17_pos N_VSSC_R17_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M22 N_VDD_M22_d N_U33_U29_c2_M22_g N_VSSC_M22_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M23 N_VDD_M22_d N_U33_U29_c2_M23_g N_VSSC_M23_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M24 N_VDD_M24_d N_U33_U29_c2_M24_g N_VSSC_M23_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_VDD_M24_d N_U33_U29_c2_M25_g N_VSSC_M25_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_VDD_M26_d N_U33_U29_c2_M26_g N_VSSC_M26_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_VDD_M26_d N_U33_U29_c2_M27_g N_VSSC_M27_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_VDD_M28_d N_U33_U29_c2_M28_g N_VSSC_M27_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_VDD_M28_d N_U33_U29_c2_M29_g N_VSSC_M22_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M3 N_VSSC_M3_d N_U34_U31_r2_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
M4 N_VSSC_M3_d N_U34_U31_r2_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M5 N_VSSC_M5_d N_U34_U31_r2_M5_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M6 N_VSSC_M5_d N_U34_U31_r2_M6_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M7 N_VSSC_M7_d N_U34_U31_r2_M7_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M8 N_VSSC_M7_d N_U34_U31_r2_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M9 N_VSSC_M9_d N_U34_U31_r2_M9_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M10 N_VSSC_M9_d N_U34_U31_r2_M10_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M11 N_VSSC_M11_d N_U34_U31_r2_M11_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M12 N_VSSC_M11_d N_U34_U31_r2_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M13 N_VSSC_M13_d N_U34_U31_r2_M13_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M14 N_VSSC_M13_d N_U34_U31_r2_M14_g N_VDD_M14_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
D30@2 N_VSSC_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSSC_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSSC_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSSC_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSSC_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSSC_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSSC_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSSC_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSSC_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC8_1 N_VDD_C8_1_pos N_U33_U29_c2_C8_1_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "pv0c.dist.sp.PV0C.pxi"
*
.ends
*
*
