* File: pc3c03.dist.sp
* Created: Sun Jul  4 12:22:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c03.dist.sp.pex"
.subckt pc3c03  CCLK VSS VDD CP VDDO VSSO
* 
M17 N_CP_M33_d N_NODE_M17_g N_VSS_M17_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M18 N_CP_M34_d N_NODE_M18_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M21 N_CP_M37_d N_NODE_M21_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M38_d N_NODE_M22_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M25 N_CP_M41_d N_NODE_M25_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M26 N_CP_M42_d N_NODE_M26_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M29 N_CP_M45_d N_NODE_M29_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M30 N_CP_M46_d N_NODE_M30_g N_VSS_M30_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M1 N_NODE_M1_d N_CCLK_M1_g N_VDD_M1_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_NODE_M1_d N_CCLK_M3_g N_VDD_M3_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M5 N_NODE_M5_d N_CCLK_M5_g N_VDD_M5_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M7 N_NODE_M5_d N_CCLK_M7_g N_VDD_M7_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M9 N_NODE_M9_d N_CCLK_M9_g N_VDD_M9_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M11 N_NODE_M9_d N_CCLK_M11_g N_VDD_M11_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M13 N_NODE_M13_d N_CCLK_M13_g N_VDD_M13_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M15 N_NODE_M13_d N_CCLK_M15_g N_VDD_M15_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M19_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M27 N_CP_M27_d N_NODE_M27_g N_VDD_M24_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M28 N_CP_M27_d N_NODE_M28_g N_VDD_M28_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M31 N_CP_M31_d N_NODE_M31_g N_VDD_M28_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M32 N_CP_M31_d N_NODE_M32_g N_VDD_M32_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M35 N_CP_M35_d N_NODE_M35_g N_VDD_M32_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M36 N_CP_M35_d N_NODE_M36_g N_VDD_M36_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M39 N_CP_M39_d N_NODE_M39_g N_VDD_M36_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M40 N_CP_M39_d N_NODE_M40_g N_VDD_M40_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M43 N_CP_M43_d N_NODE_M43_g N_VDD_M40_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M44 N_CP_M43_d N_NODE_M44_g N_VDD_M44_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M47 N_CP_M47_d N_NODE_M47_g N_VDD_M44_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M48 N_CP_M47_d N_NODE_M48_g N_VDD_M48_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D49 N_VSS_M2_b N_CCLK_D49_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M2 N_NODE_M2_d N_CCLK_M2_g N_VSS_M2_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4 N_NODE_M2_d N_CCLK_M4_g N_VSS_M4_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M33 N_CP_M33_d N_NODE_M33_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M34 N_CP_M34_d N_NODE_M34_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_NODE_M6_d N_CCLK_M6_g N_VSS_M6_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8 N_NODE_M6_d N_CCLK_M8_g N_VSS_M8_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_CP_M37_d N_NODE_M37_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M38 N_CP_M38_d N_NODE_M38_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M10 N_NODE_M10_d N_CCLK_M10_g N_VSS_M10_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M12 N_NODE_M10_d N_CCLK_M12_g N_VSS_M12_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41 N_CP_M41_d N_NODE_M41_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M42 N_CP_M42_d N_NODE_M42_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_NODE_M14_d N_CCLK_M14_g N_VSS_M14_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M16 N_NODE_M14_d N_CCLK_M16_g N_VSS_M16_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_CP_M45_d N_NODE_M45_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M46 N_CP_M46_d N_NODE_M46_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c03.dist.sp.PC3C03.pxi"
*
.ends
*
*
