* File: pv0f.dist.sp
* Created: Sun Jul  4 13:14:38 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0f.dist.sp.pex"
.subckt pv0f  VSS VDDO VDD
* 
M4 N_VDDO_M5_d N_U37_U29_c2_M4_g N_VSS_M11_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDO_M5_d N_U37_U29_c2_M5_g N_VSS_M5_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDO_M7_d N_U37_U29_c2_M6_g N_VSS_M6_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M7 N_VDDO_M7_d N_U37_U29_c2_M7_g N_VSS_M12_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDO_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U34_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U37_U29_c2_R2_pos N_noxref_6_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_6_R3_pos N_VSS_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M8 N_VDDO_M8_d N_U37_U29_c2_M8_g N_VSS_M8_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M9 N_VDDO_M8_d N_U37_U29_c2_M9_g N_VSS_M9_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M10 N_VDDO_M10_d N_U37_U29_c2_M10_g N_VSS_M9_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDO_M10_d N_U37_U29_c2_M11_g N_VSS_M11_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDO_M12_d N_U37_U29_c2_M12_g N_VSS_M12_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDO_M12_d N_U37_U29_c2_M13_g N_VSS_M13_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDO_M14_d N_U37_U29_c2_M14_g N_VSS_M13_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDO_M14_d N_U37_U29_c2_M15_g N_VSS_M8_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
dX23/D0_noxref N_VSS_X23/D0_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D1_noxref N_VSS_X23/D1_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D2_noxref N_VSS_X23/D2_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D3_noxref N_VSS_X23/D3_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D4_noxref N_VSS_X23/D4_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D5_noxref N_VSS_X23/D5_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D6_noxref N_VSS_X23/D6_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D7_noxref N_VSS_X23/D7_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D8_noxref N_VSS_X23/D8_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D9_noxref N_VSS_X23/D9_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D10_noxref N_VSS_X23/D10_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D11_noxref N_VSS_X23/D11_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D12_noxref N_VSS_X23/D12_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D13_noxref N_VSS_X23/D13_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D14_noxref N_VSS_X23/D14_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D15_noxref N_VSS_X23/D15_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D16_noxref N_VSS_X23/D16_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D17_noxref N_VSS_X23/D17_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
XC3_5 N_VDDO_C3_5_pos N_U37_U29_c2_C3_5_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSS_M16_d N_U34_U22$11_gate_M16_g N_VDDO_M16_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSS_M16_d N_U34_U22$11_gate_M17_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSS_M18_d N_U34_U22$11_gate_M18_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSS_M18_d N_U34_U22$11_gate_M19_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSS_M20_d N_U34_U22$11_gate_M20_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSS_M20_d N_U34_U22$11_gate_M21_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSS_M22_d N_U34_U22$11_gate_M22_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSS_M22_d N_U34_U22$11_gate_M23_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSS_M24_d N_U34_U22$11_gate_M24_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSS_M24_d N_U34_U22$11_gate_M25_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSS_M26_d N_U34_U22$11_gate_M26_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSS_M26_d N_U34_U22$11_gate_M27_g N_VDDO_M27_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pv0f.dist.sp.PV0F.pxi"
*
.ends
*
*
