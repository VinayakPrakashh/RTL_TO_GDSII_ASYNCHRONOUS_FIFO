* File: pc3o01hv.dist.sp
* Created: Sun Jul  4 12:37:32 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o01hv.dist.sp.pex"
.subckt pc3o01hv  PAD VSS VDDO VSSO I VDD
* 
M17 N_PAD_M23_d N_U29_U74$9_gate_M17_g N_VSSO_M17_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M24_d N_U29_U74$9_gate_M18_g N_VSSO_M18_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M19 N_PAD_M25_d N_U29_U74$9_gate_M19_g N_VSSO_M19_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U29_U74$9_gate_M20_g N_VSSO_M17_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M21 N_PAD_M15_d N_U29_U74$9_gate_M21_g N_VSSO_M21_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M22 N_PAD_M16_d N_U29_U74$9_gate_M22_g N_VSSO_M19_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR39 N_VSSO_R39_pos N_U29_U74$9_gate_R39_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR40 N_U29_U37_r2_R40_pos N_VDDO_R40_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M23 N_PAD_M23_d N_U29_U74$9_gate_M23_g N_VSSO_M23_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U29_U74$9_gate_M24_g N_VSSO_M23_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U29_U74$9_gate_M25_g N_VSSO_M25_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U29_U74$9_gate_M26_g N_VSSO_M25_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_ngate_M15_g N_VSSO_M15_s N_VSSO_M23_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_ngate_M16_g N_VSSO_M15_s N_VSSO_M23_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR13 U29_U69_padr N_noxref_2_R13_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR14 N_noxref_2_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M29 N_VDDO_M29_d N_U29_U37_r2_M29_g N_PAD_M29_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M30 N_VDDO_M31_d N_U29_U37_r2_M30_g N_PAD_M29_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M38_d N_pgate_M27_g N_PAD_M27_s N_VDDO_M31_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_pgate_M28_g N_PAD_M27_s N_VDDO_M31_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M31 N_VDDO_M31_d N_U29_U37_r2_M31_g N_PAD_M31_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U37_r2_M32_g N_PAD_M31_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U37_r2_M33_g N_PAD_M33_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U37_r2_M34_g N_PAD_M33_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_VDDO_M34_d N_U29_U37_r2_M35_g N_PAD_M35_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U29_U37_r2_M36_g N_PAD_M35_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_VDDO_M36_d N_U29_U37_r2_M37_g N_PAD_M37_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_VDDO_M38_d N_U29_U37_r2_M38_g N_PAD_M37_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M1 N_ngate_M1_d N_U28_ISHF_M1_g N_VSSO_M1_s N_VSS_M1_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M1@2 N_ngate_M1_d N_U28_ISHF_M1@2_g N_VSSO_M1@2_s N_VSS_M1_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M2 N_pgate_M2_d N_net_m2_VDDO_res_M2_g N_ngate_M2_s N_VSS_M1_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M2@2 N_pgate_M2@2_d N_net_m2_VDDO_res_M2@2_g N_ngate_M2_s N_VSS_M1_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M2@3 N_pgate_M2@2_d N_net_m2_VDDO_res_M2@3_g N_ngate_M2@3_s N_VSS_M1_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9 N_U28_U13_MPLL1_dr_M9_d N_I_M9_g N_VSSO_M9_s N_VSS_M1_b NHV L=3.6e-07
+ W=8e-06 AD=4.96e-12 AS=5.12e-12 PD=1.724e-05 PS=1.728e-05
M10 N_U28_ISHF_M10_d N_U28_U13_MPLL1_dr_M10_g N_VSSO_M10_s N_VSS_M1_b NHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M10@2 N_U28_ISHF_M10_d N_U28_U13_MPLL1_dr_M10@2_g N_VSSO_M10@2_s N_VSS_M1_b NHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@3 N_U28_ISHF_M10@3_d N_U28_U13_MPLL1_dr_M10@3_g N_VSSO_M10@2_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@4 N_U28_ISHF_M10@3_d N_U28_U13_MPLL1_dr_M10@4_g N_VSSO_M10@4_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@5 N_U28_ISHF_M10@5_d N_U28_U13_MPLL1_dr_M10@5_g N_VSSO_M10@4_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@6 N_U28_ISHF_M10@5_d N_U28_U13_MPLL1_dr_M10@6_g N_VSSO_M10@6_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M5 N_U28_U13_U6_drain_M5_d N_net_m5_VSS_res_M5_g N_VSS_M5_s N_VSS_M1_b N18
+ L=1.8e-07 W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M3 N_pgate_M3_d N_U28_ISHF_M3_g N_VDDO_M3_s N_VDDO_M3_b PHV L=3.6e-07 W=2e-05
+ AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M3@2 N_pgate_M3@2_d N_U28_ISHF_M3@2_g N_VDDO_M3_s N_VDDO_M3_b PHV L=3.6e-07
+ W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M4 N_ngate_M4_d N_net_m4_VSSO_res_M4_g N_pgate_M4_s N_VDDO_M3_b PHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4@2 N_ngate_M4_d N_net_m4_VSSO_res_M4@2_g N_pgate_M4@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M4@3 N_ngate_M4@3_d N_net_m4_VSSO_res_M4@3_g N_pgate_M4@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7 N_U28_U13_MPLL1_dr_M7_d N_I_M7_g N_VDDO_M7_s N_VDDO_M3_b PHV L=3.6e-07
+ W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M8 N_U28_ISHF_M8_d N_U28_U13_MPLL1_dr_M8_g N_VDDO_M8_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M8@2 N_U28_ISHF_M8_d N_U28_U13_MPLL1_dr_M8@2_g N_VDDO_M8@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@3 N_U28_ISHF_M8@3_d N_U28_U13_MPLL1_dr_M8@3_g N_VDDO_M8@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@4 N_U28_ISHF_M8@3_d N_U28_U13_MPLL1_dr_M8@4_g N_VDDO_M8@4_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@5 N_U28_ISHF_M8@5_d N_U28_U13_MPLL1_dr_M8@5_g N_VDDO_M8@4_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@6 N_U28_ISHF_M8@5_d N_U28_U13_MPLL1_dr_M8@6_g N_VDDO_M8@6_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M6 N_U28_U13_U6_drain_M6_d N_net_m6_VDD_res_M6_g N_VDD_M6_s N_VDD_M6_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M6@2 N_U28_U13_U6_drain_M6_d N_net_m6_VDD_res_M6@2_g N_VDD_M6@2_s N_VDD_M6_b
+ P18 L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D12 N_VSS_M1_b N_I_D12_neg DN18  AREA=1e-12 PJ=4e-06
XRM2 N_net_m2_VDDO_res_RM2_pos N_VDDO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM4 N_net_m4_VSSO_res_RM4_pos N_VSSO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM5 N_net_m5_VSS_res_RM5_pos N_VSS_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM6 N_net_m6_VDD_res_RM6_pos N_VDD_RM6_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U29_U69_padr 0 17.4974f
*
.include "pc3o01hv.dist.sp.PC3O01HV.pxi"
*
.ends
*
*
