* File: apc3d01.dist.sp
* Created: Sun Jul  4 12:03:25 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apc3d01.dist.sp.pex"
.subckt apc3d01  CIN PAD VSS AVSS AVDD AVDDO AVSSO 
* 
M7 N_CIN_M7_d N_U9_MPI1_drain_M7_g N_AVSS_M7_s N_AVSS_M7_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M15 N_PAD_M21_d N_U14_U71_r1_M15_g N_AVSSO_M15_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M22_d N_U14_U71_r1_M16_g N_AVSSO_M16_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M17 N_PAD_M23_d N_U14_U71_r1_M17_g N_AVSSO_M17_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M24_d N_U14_U71_r1_M18_g N_AVSSO_M15_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M25_d N_U14_U71_r1_M19_g N_AVSSO_M19_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M20 N_PAD_M26_d N_U14_U71_r1_M20_g N_AVSSO_M17_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR8 N_U14_U71_r1_R8_pos N_AVSSO_R8_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M21 N_PAD_M21_d N_U14_U71_r1_M21_g N_AVSSO_M21_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M22 N_PAD_M22_d N_U14_U71_r1_M22_g N_AVSSO_M21_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M23_d N_U14_U71_r1_M23_g N_AVSSO_M23_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U14_U71_r1_M24_g N_AVSSO_M23_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U14_U71_r1_M25_g N_AVSSO_M25_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U14_U71_r1_M26_g N_AVSSO_M25_s N_AVSSO_M21_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR11 N_PAD_R11_pos N_noxref_2_R11_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR12 N_noxref_2_R12_pos N_U14_padr_R12_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M27 N_AVDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M27_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M28 N_AVDDO_M31_d N_U14_pgate_tol_M28_g N_PAD_M27_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_AVDDO_M38_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_AVDDO_M30_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M31 N_AVDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_AVDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_AVDDO_M32_d N_U14_pgate_tol_M33_g N_PAD_M33_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_AVDDO_M34_d N_U14_pgate_tol_M34_g N_PAD_M33_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_AVDDO_M34_d N_U14_pgate_tol_M35_g N_PAD_M35_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_AVDDO_M36_d N_U14_pgate_tol_M36_g N_PAD_M35_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_AVDDO_M36_d N_U14_pgate_tol_M37_g N_PAD_M37_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_AVDDO_M38_d N_U14_pgate_tol_M38_g N_PAD_M37_s N_AVDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M9 N_U14_pgate_tol_M9_s N_net_m9_AVDDO_res_M9_g N_U14_pgate_tol_M9_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M9@2 N_U14_pgate_tol_M9@2_s N_net_m9_AVDDO_res_M9@2_g N_U14_pgate_tol_M9@2_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M9@3 N_U14_pgate_tol_M9@3_s N_net_m9_AVDDO_res_M9@3_g N_U14_pgate_tol_M9@3_s
+ N_AVSSO_M9_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M13 N_AVDDO_M13_d N_net_m13_AVDDO_res_M13_g N_U14_pgate_tol_M13_s N_AVSSO_M9_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M6 N_U14_padr_M6_d N_net_m6_AVSSO_res_M6_g N_AVSSO_M6_s N_AVSSO_M9_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6@2 N_U14_padr_M6@2_d N_net_m6_AVSSO_res_M6@2_g N_AVSSO_M6_s N_AVSSO_M9_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_U9_MPI1_drain_M5_d N_U14_padr_M5_g N_AVSSO_M5_s N_AVSSO_M9_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M14 N_U14_pgate_tol_M14_d N_net_m14_AVSSO_res_M14_g N_AVDDO_M14_s N_AVDDO_M14_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 N_U14_padr_M3_d N_net_m3_AVDDO_res_M3_g N_AVDDO_M3_s N_AVDDO_M14_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M1 U9_MPI2_drain N_U14_padr_M1_g N_AVDDO_M1_s N_AVDDO_M14_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M2 N_U9_MPI1_drain_M2_d N_U14_padr_M2_g U9_MPI2_drain N_AVDDO_M14_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M10 N_U14_pgate_tol_M10_s N_net_m10_AVSSO_res_M10_g N_U14_pgate_tol_M10_s
+ N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M10@2 N_U14_pgate_tol_M10@2_s N_net_m10_AVSSO_res_M10@2_g
+ N_U14_pgate_tol_M10@2_s N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M10@3 N_U14_pgate_tol_M10@3_s N_net_m10_AVSSO_res_M10@3_g
+ N_U14_pgate_tol_M10@3_s N_AVDDO_M14_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M4 N_CIN_M4_d N_U9_MPI1_drain_M4_g N_AVDD_M4_s N_AVDD_M4_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M4@2 N_CIN_M4@2_d N_U9_MPI1_drain_M4@2_g N_AVDD_M4_s N_AVDD_M4_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M4@3 N_CIN_M4@2_d N_U9_MPI1_drain_M4@3_g N_AVDD_M4@3_s N_AVDD_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M4@4 N_CIN_M4@4_d N_U9_MPI1_drain_M4@4_g N_AVDD_M4@3_s N_AVDD_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
D40@2 N_VSS_D40@2_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@3 N_VSS_D40@3_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@4 N_VSS_D40@4_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@5 N_VSS_D40@5_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@6 N_VSS_D40@6_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40@7 N_VSS_D40@7_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D40 N_VSS_D40_pos N_AVSSO_D40@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@2 N_AVSSO_D39@2_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@3 N_AVSSO_D39@3_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@4 N_AVSSO_D39@4_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@5 N_AVSSO_D39@5_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@6 N_AVSSO_D39@6_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39@7 N_AVSSO_D39@7_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D39 N_AVSSO_D39_pos N_VSS_D39@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XRM14 N_AVSSO_RM14_pos N_net_m14_AVSSO_res_RM14_neg RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM3 N_net_m3_AVDDO_res_RM3_pos N_AVDDO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM10 N_AVSSO_RM10_pos N_net_m10_AVSSO_res_RM10_neg RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM9 N_AVDDO_RM9_pos N_net_m9_AVDDO_res_RM9_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM13 N_net_m13_AVDDO_res_RM13_pos N_AVDDO_RM9_pos RPMPOLY2T w=2e-06
+ l=6.455e-06 
XRM6 N_net_m6_AVSSO_res_RM6_pos N_AVSSO_RM6_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U9_MPI2_drain 0 0.0183971f
*
.include "apc3d01.dist.sp.APC3D01.pxi"
*
.ends
*
*
* File: apv0a.dist.sp
* Created: Sun Jul  4 12:04:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apv0a.dist.sp.pex"
.subckt apv0a  AVSSO VSS AVSS AVDD AVDDO 
* 
M4 N_AVDDO_M10_d N_U31_U29_c2_M4_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_AVDDO_M11_d N_U31_U29_c2_M5_g N_AVSSO_M5_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_AVDDO_M12_d N_U31_U29_c2_M6_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_AVDDO_M13_d N_U31_U29_c2_M7_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_AVDDO_M14_d N_U31_U29_c2_M8_g N_AVSSO_M8_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_AVDDO_M15_d N_U31_U29_c2_M9_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR16 N_AVDDO_R16_pos N_noxref_3_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR17 N_noxref_3_R17_pos N_U19_U31_r2_R17_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_U31_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_AVSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_AVDDO_M10_d N_U31_U29_c2_M10_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_AVDDO_M11_d N_U31_U29_c2_M11_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_AVDDO_M12_d N_U31_U29_c2_M12_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_AVDDO_M13_d N_U31_U29_c2_M13_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_AVDDO_M14_d N_U31_U29_c2_M14_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_AVDDO_M15_d N_U31_U29_c2_M15_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M18 N_AVSSO_M18_d N_U19_U31_r2_M18_g N_AVDDO_M18_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M19 N_AVSSO_M18_d N_U19_U31_r2_M19_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_AVSSO_M20_d N_U19_U31_r2_M20_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_AVSSO_M20_d N_U19_U31_r2_M21_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_AVSSO_M22_d N_U19_U31_r2_M22_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_AVSSO_M22_d N_U19_U31_r2_M23_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_AVSSO_M24_d N_U19_U31_r2_M24_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_AVSSO_M24_d N_U19_U31_r2_M25_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_AVSSO_M26_d N_U19_U31_r2_M26_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_AVSSO_M26_d N_U19_U31_r2_M27_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M28 N_AVSSO_M28_d N_U19_U31_r2_M28_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M29 N_AVSSO_M28_d N_U19_U31_r2_M29_g N_AVDDO_M29_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
D30@2 N_AVSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_AVSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_AVSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_AVSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_AVSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_AVSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_AVSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_AVSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_AVSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC6_7 N_AVDDO_C6_7_pos N_U31_U29_c2_C6_7_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "apv0a.dist.sp.APV0A.pxi"
*
.ends
*
*
* File: apv0i.dist.sp
* Created: Sun Jul  4 12:05:08 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apv0i.dist.sp.pex"
.subckt apv0i  AVSS VSS AVDD AVDDO AVSSO 
* 
M18 N_AVDD_M24_d N_U38_U18_r1_M18_g N_AVSS_M18_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_AVDD_M25_d N_U38_U18_r1_M19_g N_AVSS_M19_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_AVDD_M26_d N_U38_U18_r1_M20_g N_AVSS_M20_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M21 N_AVDD_M27_d N_U38_U18_r1_M21_g N_AVSS_M18_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M22 N_AVDD_M28_d N_U38_U18_r1_M22_g N_AVSS_M22_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M23 N_AVDD_M29_d N_U38_U18_r1_M23_g N_AVSS_M20_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_AVDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U39_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR15 N_U38_U18_r1_R15_pos N_noxref_5_R15_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_noxref_5_R16_pos N_AVSS_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M24 N_AVDD_M24_d N_U38_U18_r1_M24_g N_AVSS_M24_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_AVDD_M25_d N_U38_U18_r1_M25_g N_AVSS_M24_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_AVDD_M26_d N_U38_U18_r1_M26_g N_AVSS_M26_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_AVDD_M27_d N_U38_U18_r1_M27_g N_AVSS_M26_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_AVDD_M28_d N_U38_U18_r1_M28_g N_AVSS_M28_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_AVDD_M29_d N_U38_U18_r1_M29_g N_AVSS_M28_s N_AVSS_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M3 N_AVSS_M3_d N_U39_U31_r2_M3_g N_AVDD_M3_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=5.68e-11 PD=4.494e-05 PS=8.284e-05
M4 N_AVSS_M3_d N_U39_U31_r2_M4_g N_AVDD_M4_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M5 N_AVSS_M5_d N_U39_U31_r2_M5_g N_AVDD_M4_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M6 N_AVSS_M5_d N_U39_U31_r2_M6_g N_AVDD_M6_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M7 N_AVSS_M7_d N_U39_U31_r2_M7_g N_AVDD_M6_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M8 N_AVSS_M7_d N_U39_U31_r2_M8_g N_AVDD_M8_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M9 N_AVSS_M9_d N_U39_U31_r2_M9_g N_AVDD_M8_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M10 N_AVSS_M9_d N_U39_U31_r2_M10_g N_AVDD_M10_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M11 N_AVSS_M11_d N_U39_U31_r2_M11_g N_AVDD_M10_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M12 N_AVSS_M11_d N_U39_U31_r2_M12_g N_AVDD_M12_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M13 N_AVSS_M13_d N_U39_U31_r2_M13_g N_AVDD_M12_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M14 N_AVSS_M13_d N_U39_U31_r2_M14_g N_AVDD_M14_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=5.68e-11 PD=4.494e-05 PS=8.284e-05
D31@2 N_AVSS_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_AVSS_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_AVSS_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_AVSS_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_AVSS_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_AVSS_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_AVSS_D31@8_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_AVSS_D31@9_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_AVSS_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@2 N_VSS_D30@2_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSS_D30@3_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSS_D30@4_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSS_D30@5_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSS_D30@6_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSS_D30@7_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSS_D30@8_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSS_D30@9_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSS_D30_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC4_10 N_AVDD_C4_10_pos N_U38_U18_r1_C4_10_neg NWCAPH2T  L=1.513e-05
+ W=1.513e-05
*
.include "apv0i.dist.sp.APV0I.pxi"
*
.ends
*
*
* File: apvda.dist.sp
* Created: Sun Jul  4 12:05:05 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apvda.dist.sp.pex"
.subckt apvda  AVDDO VSS AVSS AVDD AVSSO 
* 
M4 N_AVDDO_M10_d N_U30_U29_c2_M4_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_AVDDO_M11_d N_U30_U29_c2_M5_g N_AVSSO_M5_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_AVDDO_M12_d N_U30_U29_c2_M6_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_AVDDO_M13_d N_U30_U29_c2_M7_g N_AVSSO_M4_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_AVDDO_M14_d N_U30_U29_c2_M8_g N_AVSSO_M8_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_AVDDO_M15_d N_U30_U29_c2_M9_g N_AVSSO_M6_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR16 N_AVDDO_R16_pos N_noxref_3_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR17 N_noxref_3_R17_pos N_U19_U31_r2_R17_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_U30_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_AVSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_AVDDO_M10_d N_U30_U29_c2_M10_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_AVDDO_M11_d N_U30_U29_c2_M11_g N_AVSSO_M10_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_AVDDO_M12_d N_U30_U29_c2_M12_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_AVDDO_M13_d N_U30_U29_c2_M13_g N_AVSSO_M12_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_AVDDO_M14_d N_U30_U29_c2_M14_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_AVDDO_M15_d N_U30_U29_c2_M15_g N_AVSSO_M14_s N_AVSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M18 N_AVSSO_M18_d N_U19_U31_r2_M18_g N_AVDDO_M18_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M19 N_AVSSO_M18_d N_U19_U31_r2_M19_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_AVSSO_M20_d N_U19_U31_r2_M20_g N_AVDDO_M19_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_AVSSO_M20_d N_U19_U31_r2_M21_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_AVSSO_M22_d N_U19_U31_r2_M22_g N_AVDDO_M21_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_AVSSO_M22_d N_U19_U31_r2_M23_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_AVSSO_M24_d N_U19_U31_r2_M24_g N_AVDDO_M23_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_AVSSO_M24_d N_U19_U31_r2_M25_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_AVSSO_M26_d N_U19_U31_r2_M26_g N_AVDDO_M25_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_AVSSO_M26_d N_U19_U31_r2_M27_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M28 N_AVSSO_M28_d N_U19_U31_r2_M28_g N_AVDDO_M27_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M29 N_AVSSO_M28_d N_U19_U31_r2_M29_g N_AVDDO_M29_s N_AVDDO_M18_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
D30@2 N_AVSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_AVSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_AVSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_AVSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_AVSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_AVSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_AVSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_AVSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_AVSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_AVSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC3_7 N_AVDDO_C3_7_pos N_U30_U29_c2_C3_7_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "apvda.dist.sp.APVDA.pxi"
*
.ends
*
*
* File: apvdi.dist.sp
* Created: Sun Jul  4 12:06:27 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "apvdi.dist.sp.pex"
.subckt apvdi  AVDD VSS AVSS AVDDO AVSSO 
* 
M18 N_AVDD_M24_d N_U33_U18_r1_M18_g N_AVSSO_M18_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_AVDD_M25_d N_U33_U18_r1_M19_g N_AVSSO_M19_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_AVDD_M26_d N_U33_U18_r1_M20_g N_AVSSO_M20_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M21 N_AVDD_M27_d N_U33_U18_r1_M21_g N_AVSSO_M18_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M22 N_AVDD_M28_d N_U33_U18_r1_M22_g N_AVSSO_M22_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M23 N_AVDD_M29_d N_U33_U18_r1_M23_g N_AVSSO_M20_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_AVDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U34_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR15 N_U33_U18_r1_R15_pos N_noxref_5_R15_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_noxref_5_R16_pos N_AVSS_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M24 N_AVDD_M24_d N_U33_U18_r1_M24_g N_AVSSO_M24_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_AVDD_M25_d N_U33_U18_r1_M25_g N_AVSSO_M24_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_AVDD_M26_d N_U33_U18_r1_M26_g N_AVSSO_M26_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_AVDD_M27_d N_U33_U18_r1_M27_g N_AVSSO_M26_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_AVDD_M28_d N_U33_U18_r1_M28_g N_AVSSO_M28_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_AVDD_M29_d N_U33_U18_r1_M29_g N_AVSSO_M28_s N_AVSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
D31@2 N_AVSS_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_AVSS_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_AVSS_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_AVSS_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_AVSS_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_AVSS_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_AVSS_D31@8_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_AVSS_D31@9_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_AVSS_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@2 N_VSS_D30@2_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSS_D30@3_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSS_D30@4_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSS_D30@5_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSS_D30@6_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSS_D30@7_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSS_D30@8_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSS_D30@9_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSS_D30_pos N_AVSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC3_10 N_AVDD_C3_10_pos N_U33_U18_r1_C3_10_neg NWCAPH2T  L=1.513e-05
+ W=1.513e-05
M3 N_AVSS_M3_d N_U34_U31_r2_M3_g N_AVDD_M3_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=5.68e-11 PD=4.494e-05 PS=8.284e-05
M4 N_AVSS_M3_d N_U34_U31_r2_M4_g N_AVDD_M4_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M5 N_AVSS_M5_d N_U34_U31_r2_M5_g N_AVDD_M4_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M6 N_AVSS_M5_d N_U34_U31_r2_M6_g N_AVDD_M6_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M7 N_AVSS_M7_d N_U34_U31_r2_M7_g N_AVDD_M6_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M8 N_AVSS_M7_d N_U34_U31_r2_M8_g N_AVDD_M8_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M9 N_AVSS_M9_d N_U34_U31_r2_M9_g N_AVDD_M8_s N_AVDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M10 N_AVSS_M9_d N_U34_U31_r2_M10_g N_AVDD_M10_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M11 N_AVSS_M11_d N_U34_U31_r2_M11_g N_AVDD_M10_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M12 N_AVSS_M11_d N_U34_U31_r2_M12_g N_AVDD_M12_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M13 N_AVSS_M13_d N_U34_U31_r2_M13_g N_AVDD_M12_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=3.64e-11 PD=4.494e-05 PS=4.182e-05
M14 N_AVSS_M13_d N_U34_U31_r2_M14_g N_AVDD_M14_s N_AVDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=9.88e-11 AS=5.68e-11 PD=4.494e-05 PS=8.284e-05
*
.include "apvdi.dist.sp.APVDI.pxi"
*
.ends
*
*
* File: pc3b01d.dist.sp
* Created: Sun Jul  4 12:08:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b01d.dist.sp.pex"
.subckt pc3b01d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M56 N_U27_padr_M56_d N_net_m56_VDDO_res_M56_g U28_U22_source N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M57 U28_U22_source N_net_m57_VDDO_res_M57_g N_VSSO_M57_s N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM56 N_net_m56_VDDO_res_RM56_pos N_VDDO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM57 N_VDDO_RM56_neg N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M63 N_U27_padr_M63_d N_net_m63_VSSO_res_M63_g N_VSSO_M63_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M63@2 N_U27_padr_M63@2_d N_net_m63_VSSO_res_M63@2_g N_VSSO_M63_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62 N_U26_MPI1_drain_M62_d N_U27_padr_M62_g N_VSSO_M62_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M64 N_CIN_M64_d N_U26_MPI1_drain_M64_g N_VSS_M64_s N_VSS_M25_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M60 N_U27_padr_M60_d N_net_m60_VDDO_res_M60_g N_VDDO_M60_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 U26_MPI2_drain N_U27_padr_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M59 N_U26_MPI1_drain_M59_d N_U27_padr_M59_g U26_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M61 N_CIN_M61_d N_U26_MPI1_drain_M61_g N_VDD_M61_s N_VDD_M42_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M61@2 N_CIN_M61@2_d N_U26_MPI1_drain_M61@2_g N_VDD_M61_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M61@3 N_CIN_M61@2_d N_U26_MPI1_drain_M61@3_g N_VDD_M61@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M61@4 N_CIN_M61@4_d N_U26_MPI1_drain_M61@4_g N_VDD_M61@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM60 N_net_m60_VDDO_res_RM60_pos N_VDDO_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b01d.dist.sp.PC3B01D.pxi"
*
.ends
*
*
* File: pc3b01.dist.sp
* Created: Sun Jul  4 12:06:31 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b01.dist.sp.pex"
.subckt pc3b01  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M61 N_U27_padr_M61_d N_net_m61_VSSO_res_M61_g N_VSSO_M61_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M61@2 N_U27_padr_M61@2_d N_net_m61_VSSO_res_M61@2_g N_VSSO_M61_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60 N_U26_MPI1_drain_M60_d N_U27_padr_M60_g N_VSSO_M60_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M62 N_CIN_M62_d N_U26_MPI1_drain_M62_g N_VSS_M62_s N_VSS_M25_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 N_U27_padr_M58_d N_net_m58_VDDO_res_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M56 U26_MPI2_drain N_U27_padr_M56_g N_VDDO_M56_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M57 N_U26_MPI1_drain_M57_d N_U27_padr_M57_g U26_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M59 N_CIN_M59_d N_U26_MPI1_drain_M59_g N_VDD_M59_s N_VDD_M42_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M59@2 N_CIN_M59@2_d N_U26_MPI1_drain_M59@2_g N_VDD_M59_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M59@3 N_CIN_M59@2_d N_U26_MPI1_drain_M59@3_g N_VDD_M59@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M59@4 N_CIN_M59@4_d N_U26_MPI1_drain_M59@4_g N_VDD_M59@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM58 N_net_m58_VDDO_res_RM58_pos N_VDDO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM61 N_VSSO_RM61_pos N_net_m61_VSSO_res_RM61_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b01.dist.sp.PC3B01.pxi"
*
.ends
*
*
* File: pc3b01u.dist.sp
* Created: Sun Jul  4 12:08:11 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b01u.dist.sp.pex"
.subckt pc3b01u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M35 N_PAD_M36_d N_U27_U69$9_gate_M35_g N_VSSO_M35_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U27_U69$9_gate_M36_g N_VSSO_M36_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M37 N_PAD_M38_d N_U27_U69$9_gate_M37_g N_VSSO_M37_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M38_d N_U27_U69$9_gate_M38_g N_VSSO_M35_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M39 N_PAD_M40_d N_U27_U69$9_gate_M39_g N_VSSO_M39_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U27_U69$9_gate_M40_g N_VSSO_M37_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M42_d N_U27_U69$9_gate_M41_g N_VSSO_M41_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M42_d N_U27_U69$9_gate_M42_g N_VSSO_M39_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M43_d N_U15_ngate_M33_g N_VSSO_M33_s N_VSSO_M36_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M43 N_PAD_M43_d N_U27_U69$9_gate_M43_g N_VSSO_M41_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M44 N_PAD_M34_d N_U27_U69$9_gate_M44_g N_VSSO_M44_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M34_d N_U15_ngate_M34_g N_VSSO_M33_s N_VSSO_M36_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U27_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M63_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M58 N_U15_pgate_M58_d N_net_m58_VSSO_res_M58_g N_U27_U72_pgate_M58_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M58@2 N_U15_pgate_M58_d N_net_m58_VSSO_res_M58@2_g N_U27_U72_pgate_M58@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@3 N_U15_pgate_M58@3_d N_net_m58_VSSO_res_M58@3_g N_U27_U72_pgate_M58@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@4 N_U15_pgate_M58@3_d N_net_m58_VSSO_res_M58@4_g N_U27_U72_pgate_M58@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@5 N_U15_pgate_M58@5_d N_net_m58_VSSO_res_M58@5_g N_U27_U72_pgate_M58@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U27_U69$9_gate_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XR59 N_noxref_2_R59_pos N_PAD_R59_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR60 N_noxref_2_R60_pos N_U27_padr_R60_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M47 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M47_g N_PAD_M47_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M48 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M48_g N_PAD_M47_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M45 N_VDDO_M56_d N_U27_U72_pgate_M45_g N_PAD_M45_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M46 N_VDDO_M46_d N_U27_U72_pgate_M46_g N_PAD_M45_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M49 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M49_g N_PAD_M49_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M50_g N_PAD_M49_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M51 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M51_g N_PAD_M51_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M52_g N_PAD_M51_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M53_g N_PAD_M53_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U27_U71_UN_P_TOP_M54_g N_PAD_M53_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_VDDO_M54_d N_U27_U71_UN_P_TOP_M55_g N_PAD_M55_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M56 N_VDDO_M56_d N_U27_U71_UN_P_TOP_M56_g N_PAD_M55_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M57 N_U15_pgate_M57_d N_net_m57_VDDO_res_M57_g N_U27_U72_pgate_M57_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M57@2 N_U15_pgate_M57_d N_net_m57_VDDO_res_M57@2_g N_U27_U72_pgate_M57@2_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M57@3 N_U15_pgate_M57@3_d N_net_m57_VDDO_res_M57@3_g N_U27_U72_pgate_M57@2_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U27_U71_UN_P_TOP_M62_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_U27_padr_M7_d N_net_m7_VSSO_res_M7_g N_VSSO_M7_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7@2 N_U27_padr_M7@2_d N_net_m7_VSSO_res_M7@2_g N_VSSO_M7_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6 N_U26_MPI1_drain_M6_d N_U27_padr_M6_g N_VSSO_M6_s N_VSS_M57_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M8 N_CIN_M8_d N_U26_MPI1_drain_M8_g N_VSS_M8_s N_VSS_M57_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M30 N_U15_U12_oenb_M30_d N_U15_U15_OUTSHIFT_M30_g N_VSSO_M30_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M9 N_U15_ngate_M9_d N_U15_ISHF_M9_g N_VSSO_M9_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9@2 N_U15_ngate_M9_d N_U15_ISHF_M9@2_g N_VSSO_M9@2_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M29 N_U15_ngate_M29_d N_U15_U15_OUTSHIFT_M29_g N_VSSO_M9@2_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M10 N_U15_pgate_M10_d N_U15_U12_oenb_M10_g N_U15_ngate_M10_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M10@2 N_U15_pgate_M10@2_d N_U15_U12_oenb_M10@2_g N_U15_ngate_M10_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M10@3 N_U15_pgate_M10@2_d N_U15_U12_oenb_M10@3_g N_U15_ngate_M10@3_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M23 N_U15_U15_MPLL1_dr_M23_d N_OEN_M23_g N_VSSO_M23_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M25 N_VDDO_M25_d N_U15_U15_MN1_drai_M25_g N_U15_U15_MPLL1_dr_M25_s N_VSS_M57_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M23@2 N_U15_U15_MPLL1_dr_M23@2_d N_OEN_M23@2_g N_VSSO_M23_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M24 N_U15_U15_OUTSHIFT_M24_d N_U15_U15_MN1_drai_M24_g N_VSSO_M24_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M24@2 N_U15_U15_OUTSHIFT_M24@2_d N_U15_U15_MN1_drai_M24@2_g N_VSSO_M24_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M17 N_VDDO_M17_d N_U15_U14_MN1_drai_M17_g N_U15_U14_MPLL1_dr_M17_s N_VSS_M57_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M15 N_U15_U14_MPLL1_dr_M15_d N_I_M15_g N_VSSO_M15_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M15@2 N_U15_U14_MPLL1_dr_M15@2_d N_I_M15@2_g N_VSSO_M15_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U15_ISHF_M16_d N_U15_U14_MN1_drai_M16_g N_VSSO_M16_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16@2 N_U15_ISHF_M16@2_d N_U15_U14_MN1_drai_M16@2_g N_VSSO_M16_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M18 N_U15_U14_MN1_drai_M18_d N_I_M18_g N_VSS_M18_s N_VSS_M57_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M26 N_U15_U15_MN1_drai_M26_d N_OEN_M26_g N_VSS_M18_s N_VSS_M57_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U27_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M4 N_U27_padr_M4_d N_net_m4_VDDO_res_M4_g N_VDDO_M4_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M2 U26_MPI2_drain N_U27_padr_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M3 N_U26_MPI1_drain_M3_d N_U27_padr_M3_g U26_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M31 N_U15_U12_oenb_M31_d N_U15_U15_OUTSHIFT_M31_g N_VDDO_M31_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M31@2 N_U15_U12_oenb_M31@2_d N_U15_U15_OUTSHIFT_M31@2_g N_VDDO_M31_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M11 N_U15_pgate_M11_d N_U15_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M11@2 N_U15_pgate_M11@2_d N_U15_ISHF_M11@2_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M32 N_U15_pgate_M11@2_d N_U15_U12_oenb_M32_g N_VDDO_M32_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M32@2 N_U15_pgate_M32@2_d N_U15_U12_oenb_M32@2_g N_VDDO_M32_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M12 N_U15_ngate_M12_d N_U15_U15_OUTSHIFT_M12_g N_U15_pgate_M12_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M12@2 N_U15_ngate_M12_d N_U15_U15_OUTSHIFT_M12@2_g N_U15_pgate_M12@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M12@3 N_U15_ngate_M12@3_d N_U15_U15_OUTSHIFT_M12@3_g N_U15_pgate_M12@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M21 N_U15_U15_MPLL1_dr_M21_d N_U15_U15_OUTSHIFT_M21_g N_VDDO_M21_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M22 N_U15_U15_OUTSHIFT_M22_d N_U15_U15_MPLL1_dr_M22_g N_VDDO_M21_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M13 N_U15_U14_MPLL1_dr_M13_d N_U15_ISHF_M13_g N_VDDO_M13_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M14 N_U15_ISHF_M14_d N_U15_U14_MPLL1_dr_M14_g N_VDDO_M13_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M5 N_CIN_M5_d N_U26_MPI1_drain_M5_g N_VDD_M5_s N_VDD_M19_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M5@2 N_CIN_M5@2_d N_U26_MPI1_drain_M5@2_g N_VDD_M5_s N_VDD_M19_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M5@3 N_CIN_M5@2_d N_U26_MPI1_drain_M5@3_g N_VDD_M5@3_s N_VDD_M19_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M5@4 N_CIN_M5@4_d N_U26_MPI1_drain_M5@4_g N_VDD_M5@3_s N_VDD_M19_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M19 N_U15_U14_MN1_drai_M19_d N_I_M19_g N_VDD_M19_s N_VDD_M19_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M19@2 N_U15_U14_MN1_drai_M19_d N_I_M19@2_g N_VDD_M19@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M27 N_U15_U15_MN1_drai_M27_d N_OEN_M27_g N_VDD_M19@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M27@2 N_U15_U15_MN1_drai_M27_d N_OEN_M27@2_g N_VDD_M27@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D20 N_VSS_M57_b N_I_D20_neg DN18  AREA=2.5e-13 PJ=2e-06
D28 N_VSS_M57_b N_OEN_D28_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_net_m4_VDDO_res_RM4_pos N_VDDO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM57 N_VDDO_RM57_pos N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM7 N_VSSO_RM7_pos N_net_m7_VSSO_res_RM7_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM58 N_net_m58_VSSO_res_RM58_pos N_VSSO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b01u.dist.sp.PC3B01U.pxi"
*
.ends
*
*
* File: pc3b02d.dist.sp
* Created: Sun Jul  4 12:09:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b02d.dist.sp.pex"
.subckt pc3b02d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M69 N_U27_padr_M69_d N_net_m69_VDDO_res_M69_g U28_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U28_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U27_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U27_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U26_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M68 N_CIN_M68_d N_U26_MPI1_drain_M68_g N_VSS_M68_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U26_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U26_MPI1_drain_M63_d N_U27_padr_M63_g U26_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M65 N_CIN_M65_d N_U26_MPI1_drain_M65_g N_VDD_M65_s N_VDD_M48_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M65@2 N_CIN_M65@2_d N_U26_MPI1_drain_M65@2_g N_VDD_M65_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@3 N_CIN_M65@2_d N_U26_MPI1_drain_M65@3_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@4 N_CIN_M65@4_d N_U26_MPI1_drain_M65@4_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.360765f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b02d.dist.sp.PC3B02D.pxi"
*
.ends
*
*
* File: pc3b02.dist.sp
* Created: Sun Jul  4 12:09:55 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b02.dist.sp.pex"
.subckt pc3b02  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U27_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U27_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U26_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M68 N_CIN_M68_d N_U26_MPI1_drain_M68_g N_VSS_M68_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U26_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U26_MPI1_drain_M63_d N_U27_padr_M63_g U26_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M65 N_CIN_M65_d N_U26_MPI1_drain_M65_g N_VDD_M65_s N_VDD_M48_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M65@2 N_CIN_M65@2_d N_U26_MPI1_drain_M65@2_g N_VDD_M65_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@3 N_CIN_M65@2_d N_U26_MPI1_drain_M65@3_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@4 N_CIN_M65@4_d N_U26_MPI1_drain_M65@4_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.360765f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b02.dist.sp.PC3B02.pxi"
*
.ends
*
*
* File: pc3b02u.dist.sp
* Created: Sun Jul  4 12:11:25 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b02u.dist.sp.pex"
.subckt pc3b02u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M69 N_U27_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M37_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VSSO_res_RM69_pos N_VSSO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U27_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U27_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U26_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M68 N_CIN_M68_d N_U26_MPI1_drain_M68_g N_VSS_M68_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U26_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U26_MPI1_drain_M63_d N_U27_padr_M63_g U26_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M65 N_CIN_M65_d N_U26_MPI1_drain_M65_g N_VDD_M65_s N_VDD_M48_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M65@2 N_CIN_M65@2_d N_U26_MPI1_drain_M65@2_g N_VDD_M65_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@3 N_CIN_M65@2_d N_U26_MPI1_drain_M65@3_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M65@4 N_CIN_M65@4_d N_U26_MPI1_drain_M65@4_g N_VDD_M65@3_s N_VDD_M48_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.360765f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b02u.dist.sp.PC3B02U.pxi"
*
.ends
*
*
* File: pc3b03d.dist.sp
* Created: Sun Jul  4 12:13:10 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b03d.dist.sp.pex"
.subckt pc3b03d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M71 N_U28_padr_M71_d N_net_m71_VDDO_res_M71_g U29_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U29_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b03d.dist.sp.PC3B03D.pxi"
*
.ends
*
*
* File: pc3b03ed.dist.sp
* Created: Sun Jul  4 12:13:05 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b03ed.dist.sp.pex"
.subckt pc3b03ed  PAD I OEN CIN RENB VDD VSS VDDO VSSO 
* 
M81 U30_U22_source N_U30_MN3_drain_M81_g N_VSSO_M81_s N_VSS_M31_b NHV L=5.5e-06
+ W=1.33e-06 AD=2.66e-13 AS=1.0374e-12 PD=1.73e-06 PS=4.22e-06
M71 N_U30_MN3_drain_M71_d N_U30_U24_OUTSHIFT_M71_g N_VSSO_M71_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M80 N_U28_padr_M80_d N_U30_MN3_drain_M80_g U30_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=1.33e-06 AD=1.0374e-12 AS=2.66e-13 PD=4.22e-06 PS=1.73e-06
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M72 N_U30_MN3_drain_M72_d N_U30_U24_OUTSHIFT_M72_g N_VDDO_M72_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M75 N_U30_U24_OUTSHIFT_M75_d N_U30_U24_U6_drain_M75_g N_VDDO_M75_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
M74 N_U30_U24_U6_drain_M74_d N_U30_U24_OUTSHIFT_M74_g N_VDDO_M75_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_4_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_4_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_RM31_neg N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M77 N_U30_U24_OUTSHIFT_M77_d N_U30_U24_nsgate_M77_g N_VSSO_M77_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M76 N_U30_U24_U6_drain_M76_d N_RENB_M76_g N_VSSO_M76_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M73 N_U30_U24_nsgate_M73_d N_RENB_M73_g N_VSS_M73_s N_VSS_M31_b N18 L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M78_b PHV L=3.6e-07
+ W=8.06e-06 AD=5.4002e-12 AS=3.3046e-12 PD=1.746e-05 PS=8.88e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M78_b PHV
+ L=3.6e-07 W=8.06e-06 AD=3.3046e-12 AS=3.3046e-12 PD=8.88e-06 PS=8.88e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M78_b PHV
+ L=3.6e-07 W=8.06e-06 AD=3.3046e-12 AS=3.3046e-12 PD=8.88e-06 PS=8.88e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M78_b PHV
+ L=3.6e-07 W=8.06e-06 AD=4.9972e-12 AS=3.3046e-12 PD=1.736e-05 PS=8.88e-06
M78 N_U30_U24_nsgate_M78_d N_RENB_M78_g N_VDD_M78_s N_VDD_M78_b P18 L=2e-07
+ W=2.78e-06 AD=1.946e-12 AS=1.946e-12 PD=6.96e-06 PS=6.96e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M78_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M78_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M78_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M78_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D79 N_VSS_M31_b N_RENB_D79_neg DN18  AREA=1e-12 PJ=4e-06
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U30_U22_source 0 0.0178743f
c_2 U17_U15_U8_sourc 0 0.359728f
c_3 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b03ed.dist.sp.PC3B03ED.pxi"
*
.ends
*
*
* File: pc3b03.dist.sp
* Created: Sun Jul  4 12:11:35 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b03.dist.sp.pex"
.subckt pc3b03  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b03.dist.sp.PC3B03.pxi"
*
.ends
*
*
* File: pc3b03u.dist.sp
* Created: Sun Jul  4 12:14:42 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b03u.dist.sp.pex"
.subckt pc3b03u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M71 N_U28_padr_M71_d N_net_m71_VSSO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VSSO_res_RM71_pos N_VSSO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b03u.dist.sp.PC3B03U.pxi"
*
.ends
*
*
* File: pc3b04d.dist.sp
* Created: Sun Jul  4 12:16:32 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b04d.dist.sp.pex"
.subckt pc3b04d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M71 N_U28_padr_M71_d N_net_m71_VDDO_res_M71_g U30_U22_source N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U30_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X36/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X36/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b04d.dist.sp.PC3B04D.pxi"
*
.ends
*
*
* File: pc3b04.dist.sp
* Created: Sun Jul  4 12:14:44 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b04.dist.sp.pex"
.subckt pc3b04  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X32/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X32/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b04.dist.sp.PC3B04.pxi"
*
.ends
*
*
* File: pc3b04u.dist.sp
* Created: Sun Jul  4 12:16:19 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b04u.dist.sp.pex"
.subckt pc3b04u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M71 N_U28_padr_M71_d N_net_m71_VSSO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VSSO_res_RM71_pos N_VSSO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X34/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X34/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b04u.dist.sp.PC3B04U.pxi"
*
.ends
*
*
* File: pc3b05d.dist.sp
* Created: Sun Jul  4 12:18:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b05d.dist.sp.pex"
.subckt pc3b05d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M71 N_U29_padr_M71_d N_net_m71_VDDO_res_M71_g U31_U22_source N_VSS_M43_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U31_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M43_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M39 N_PAD_M37_d N_U30_ngate_M39_g N_VSSO_M39_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M37 N_PAD_M37_d N_U29_U42_r1_M37_g N_VSSO_M37_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M40 N_PAD_M41_d N_U30_ngate_M40_g N_VSSO_M40_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M41_d N_U30_ngate_M41_g N_VSSO_M39_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M42_d N_U17_ngate2_M33_g N_VSSO_M33_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M42_d N_U30_ngate_M42_g N_VSSO_M40_s N_VSSO_M37_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M34 N_PAD_M35_d N_U17_ngate2_M34_g N_VSSO_M34_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M35_d N_U17_ngate2_M35_g N_VSSO_M33_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M31 N_PAD_M36_d N_U29_ngate3_M31_g N_VSSO_M31_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U17_ngate2_M36_g N_VSSO_M34_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M32_d N_U29_U42_r1_M38_g N_VSSO_M38_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M32 N_PAD_M32_d N_U29_ngate3_M32_g N_VSSO_M31_s N_VSSO_M37_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M44 N_U30_pgate_M44_d N_net_m44_VSSO_res_M44_g N_U29_U72_pgate_M44_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M44@2 N_U30_pgate_M44_d N_net_m44_VSSO_res_M44@2_g N_U29_U72_pgate_M44@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@3 N_U30_pgate_M44@3_d N_net_m44_VSSO_res_M44@3_g N_U29_U72_pgate_M44@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@4 N_U30_pgate_M44@3_d N_net_m44_VSSO_res_M44@4_g N_U29_U72_pgate_M44@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M44@5 N_U30_pgate_M44@5_d N_net_m44_VSSO_res_M44@5_g N_U29_U72_pgate_M44@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U29_U42_r1_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR45 N_noxref_2_R45_pos N_PAD_R45_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR46 N_noxref_2_R46_pos N_U29_padr_R46_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M59 N_VDDO_M59_d N_U29_U71_UN_P_TOP_M59_g N_PAD_M59_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M60 N_VDDO_M51_d N_U29_U71_UN_P_TOP_M60_g N_PAD_M59_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M49 N_VDDO_M58_d N_U29_U72_pgate_M49_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M50_d N_U29_U72_pgate_M50_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M51 N_VDDO_M51_d N_U29_U72_pgate_M51_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U29_U72_pgate_M52_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U29_U72_pgate_M53_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U29_U72_pgate_M54_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_VDDO_M54_d N_U29_U72_pgate_M55_g N_PAD_M55_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M56 N_VDDO_M56_d N_U29_U72_pgate_M56_g N_PAD_M55_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M57 N_VDDO_M56_d N_U29_U72_pgate_M57_g N_PAD_M57_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M58 N_VDDO_M58_d N_U29_U72_pgate_M58_g N_PAD_M57_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_U30_pgate_M43_d N_net_m43_VDDO_res_M43_g N_U29_U72_pgate_M43_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M43@2 N_U30_pgate_M43_d N_net_m43_VDDO_res_M43@2_g N_U29_U72_pgate_M43@2_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M43@3 N_U30_pgate_M43@3_d N_net_m43_VDDO_res_M43@3_g N_U29_U72_pgate_M43@2_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U29_U71_UN_P_TOP_M62_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M43_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M48 N_U29_ngate3_M48_d N_U17_ngatex_M48_g N_VSSO_M48_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M43_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M43_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M28 N_U30_U12_oenb_M28_d N_U30_U15_OUTSHIFT_M28_g N_VSSO_M28_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M9 N_U30_ngate_M9_d N_U30_ISHF_M9_g N_VSSO_M9_s N_VSS_M43_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M9@2 N_U30_ngate_M9_d N_U30_ISHF_M9@2_g N_VSSO_M9@2_s N_VSS_M43_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M27 N_U30_ngate_M27_d N_U30_U15_OUTSHIFT_M27_g N_VSSO_M9@2_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M10 N_U30_pgate_M10_d N_U30_U12_oenb_M10_g N_U30_ngate_M10_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M10@2 N_U30_pgate_M10@2_d N_U30_U12_oenb_M10@2_g N_U30_ngate_M10_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M10@3 N_U30_pgate_M10@2_d N_U30_U12_oenb_M10@3_g N_U30_ngate_M10@3_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M21 N_U30_U15_MPLL1_dr_M21_d N_OEN_M21_g N_VSSO_M21_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M23 N_VDDO_M23_d N_U30_U15_MN1_drai_M23_g N_U30_U15_MPLL1_dr_M23_s N_VSS_M43_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M21@2 N_U30_U15_MPLL1_dr_M21@2_d N_OEN_M21@2_g N_VSSO_M21_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22 N_U30_U15_OUTSHIFT_M22_d N_U30_U15_MN1_drai_M22_g N_VSSO_M22_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22@2 N_U30_U15_OUTSHIFT_M22@2_d N_U30_U15_MN1_drai_M22@2_g N_VSSO_M22_s
+ N_VSS_M43_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M15 N_VDDO_M15_d N_U30_U14_MN1_drai_M15_g N_U30_U14_MPLL1_dr_M15_s N_VSS_M43_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U30_U14_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M43_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U30_U14_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U30_ISHF_M14_d N_U30_U14_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M43_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U30_ISHF_M14@2_d N_U30_U14_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M43_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U30_U14_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M43_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M24 N_U30_U15_MN1_drai_M24_d N_OEN_M24_g N_VSS_M16_s N_VSS_M43_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U29_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M63_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M63_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M47 N_U29_ngate3_M47_d N_U17_ngatex_M47_g N_U17_ngate2_M47_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M29 N_U30_U12_oenb_M29_d N_U30_U15_OUTSHIFT_M29_g N_VDDO_M29_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M29@2 N_U30_U12_oenb_M29@2_d N_U30_U15_OUTSHIFT_M29@2_g N_VDDO_M29_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M7 N_U30_pgate_M7_d N_U30_ISHF_M7_g N_VDDO_M7_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M7@2 N_U30_pgate_M7_d N_U30_ISHF_M7@2_g N_VDDO_M7@2_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M7@3 N_U30_pgate_M7@3_d N_U30_ISHF_M7@3_g N_VDDO_M7@2_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M30 N_U30_pgate_M7@3_d N_U30_U12_oenb_M30_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M30@2 N_U30_pgate_M30@2_d N_U30_U12_oenb_M30@2_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8 N_U30_ngate_M8_d N_U30_U15_OUTSHIFT_M8_g N_U30_pgate_M8_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8@2 N_U30_ngate_M8_d N_U30_U15_OUTSHIFT_M8@2_g N_U30_pgate_M8@2_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_U30_ngate_M8@3_d N_U30_U15_OUTSHIFT_M8@3_g N_U30_pgate_M8@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M19 N_U30_U15_MPLL1_dr_M19_d N_U30_U15_OUTSHIFT_M19_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M20 N_U30_U15_OUTSHIFT_M20_d N_U30_U15_MPLL1_dr_M20_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U30_U14_MPLL1_dr_M11_d N_U30_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U30_ISHF_M12_d N_U30_U14_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M17_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M17_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M17 N_U30_U14_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U30_U14_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25 N_U30_U15_MN1_drai_M25_d N_OEN_M25_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25@2 N_U30_U15_MN1_drai_M25_d N_OEN_M25@2_g N_VDD_M25@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D18 N_VSS_M43_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
D26 N_VSS_M43_b N_OEN_D26_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM43 N_VDDO_RM43_pos N_net_m43_VDDO_res_RM43_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM44 N_net_m44_VSSO_res_RM44_pos N_VSSO_RM44_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b05d.dist.sp.PC3B05D.pxi"
*
.ends
*
*
* File: pc3b05.dist.sp
* Created: Sun Jul  4 12:17:49 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b05.dist.sp.pex"
.subckt pc3b05  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b05.dist.sp.PC3B05.pxi"
*
.ends
*
*
* File: pc3b05u.dist.sp
* Created: Sun Jul  4 12:19:24 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b05u.dist.sp.pex"
.subckt pc3b05u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M71 N_U29_padr_M71_d N_net_m71_VSSO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_VSSO_RM71_pos N_net_m71_VSSO_res_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pc3b05u.dist.sp.PC3B05U.pxi"
*
.ends
*
*
* File: pc3b21eu.dist.sp
* Created: Sun Jul  4 12:19:28 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b21eu.dist.sp.pex"
.subckt pc3b21eu  PAD I OEN RENB CIN VDD VSS VDDO VSSO 
* 
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M73 N_U27_padr_M73_d N_U32_U1_OUTSHIFT_M73_g N_VDDO_M73_s N_VDDO_M31_b PHV
+ L=2e-06 W=2e-06 AD=4.26e-12 AS=4.24e-12 PD=8.26e-06 PS=8.24e-06
M68 N_U32_U1_OUTSHIFT_M68_d N_U32_U1_U6_drain_M68_g N_VDDO_M68_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
M67 N_U32_U1_U6_drain_M67_d N_U32_U1_OUTSHIFT_M67_g N_VDDO_M68_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M58 N_U27_padr_M58_d N_net_m58_VSSO_res_M58_g N_VSSO_M58_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M58@2 N_U27_padr_M58@2_d N_net_m58_VSSO_res_M58@2_g N_VSSO_M58_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M57 N_U26_U36_drain_M57_d N_U27_padr_M57_g N_U26_U34_drain_M57_s N_VSS_M25_b
+ NHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M60 N_CIN_M60_d N_U26_U36_drain_M60_g N_VSS_M60_s N_VSS_M25_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M59 N_VDDO_M59_d N_U26_U36_drain_M59_g N_U26_U34_drain_M59_s N_VSS_M25_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M56 N_U26_U34_drain_M56_d N_U27_padr_M56_g N_VSSO_M56_s N_VSS_M25_b NHV
+ L=3.6e-07 W=9.5e-06 AD=5.89e-12 AS=5.89e-12 PD=2.024e-05 PS=2.024e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M70 N_U32_U1_OUTSHIFT_M70_d N_U32_U1_nsgate_M70_g N_VSSO_M70_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U32_U1_U6_drain_M69_d N_RENB_M69_g N_VSSO_M69_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M66 N_U32_U1_nsgate_M66_d N_RENB_M66_g N_VSS_M66_s N_VSS_M25_b N18 L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M63 N_U27_padr_M63_d N_net_m63_VDDO_res_M63_g N_VDDO_M63_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 N_U26_U30_source_M62_d N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=8.8e-12 PD=1.182e-05 PS=2.36e-05
M61 N_U26_U36_drain_M61_d N_U27_padr_M61_g N_U26_U30_source_M62_d N_VDDO_M31_b
+ PHV L=3.6e-07 W=1.1e-05 AD=6.93e-12 AS=4.51e-12 PD=2.326e-05 PS=1.182e-05
M64 N_VSSO_M64_d N_U26_U36_drain_M64_g N_U26_U30_source_M64_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M65 N_CIN_M65_d N_U26_U36_drain_M65_g N_VDD_M65_s N_VDD_M71_b PHV L=3.6e-07
+ W=9e-06 AD=6.03e-12 AS=3.69e-12 PD=1.934e-05 PS=9.82e-06
M65@2 N_CIN_M65@2_d N_U26_U36_drain_M65@2_g N_VDD_M65_s N_VDD_M71_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M65@3 N_CIN_M65@2_d N_U26_U36_drain_M65@3_g N_VDD_M65@3_s N_VDD_M71_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M65@4 N_CIN_M65@4_d N_U26_U36_drain_M65@4_g N_VDD_M65@3_s N_VDD_M71_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M71 N_U32_U1_nsgate_M71_d N_RENB_M71_g N_VDD_M71_s N_VDD_M71_b P18 L=2e-07
+ W=2.78e-06 AD=1.946e-12 AS=1.946e-12 PD=6.96e-06 PS=6.96e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M71_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M71_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M71_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M71_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D72 N_VSS_M25_b N_RENB_D72_neg DN18  AREA=1e-12 PJ=4e-06
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM63 N_net_m63_VDDO_res_RM63_pos N_VDDO_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM58 N_VSSO_RM58_pos N_net_m58_VSSO_res_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3b21eu.dist.sp.PC3B21EU.pxi"
*
.ends
*
*
* File: pc3b25eu.dist.sp
* Created: Sun Jul  4 12:21:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3b25eu.dist.sp.pex"
.subckt pc3b25eu  I OEN CIN RENB PAD VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M81 N_U29_padr_M81_d N_U32_U1_OUTSHIFT_M81_g N_VDDO_M81_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4.26e-12 AS=4.24e-12 PD=8.26e-06 PS=8.24e-06
M76 N_U32_U1_OUTSHIFT_M76_d N_U32_U1_U6_drain_M76_g N_VDDO_M76_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
M75 N_U32_U1_U6_drain_M75_d N_U32_U1_OUTSHIFT_M75_g N_VDDO_M76_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M66 N_U29_padr_M66_d N_net_m66_VSSO_res_M66_g N_VSSO_M66_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66@2 N_U29_padr_M66@2_d N_net_m66_VSSO_res_M66@2_g N_VSSO_M66_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M65 N_U26_U36_drain_M65_d N_U29_padr_M65_g N_U26_U34_drain_M65_s N_VSS_M19_b
+ NHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M68 N_CIN_M68_d N_U26_U36_drain_M68_g N_VSS_M68_s N_VSS_M19_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_VDDO_M67_d N_U26_U36_drain_M67_g N_U26_U34_drain_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M64 N_U26_U34_drain_M64_d N_U29_padr_M64_g N_VSSO_M64_s N_VSS_M19_b NHV
+ L=3.6e-07 W=9.5e-06 AD=5.89e-12 AS=5.89e-12 PD=2.024e-05 PS=2.024e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M78 N_U32_U1_OUTSHIFT_M78_d N_U32_U1_nsgate_M78_g N_VSSO_M78_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M77 N_U32_U1_U6_drain_M77_d N_RENB_M77_g N_VSSO_M77_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M74 N_U32_U1_nsgate_M74_d N_RENB_M74_g N_VSS_M74_s N_VSS_M19_b N18 L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.9e-12 PD=1.116e-05 PS=5.76e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M71 N_U29_padr_M71_d N_net_m71_VDDO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M70 N_U26_U30_source_M70_d N_U29_padr_M70_g N_VDDO_M70_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=8.8e-12 PD=1.182e-05 PS=2.36e-05
M69 N_U26_U36_drain_M69_d N_U29_padr_M69_g N_U26_U30_source_M70_d N_VDDO_M39_b
+ PHV L=3.6e-07 W=1.1e-05 AD=6.93e-12 AS=4.51e-12 PD=2.326e-05 PS=1.182e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M72 N_VSSO_M72_d N_U26_U36_drain_M72_g N_U26_U30_source_M72_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M73 N_CIN_M73_d N_U26_U36_drain_M73_g N_VDD_M73_s N_VDD_M79_b PHV L=3.6e-07
+ W=9e-06 AD=6.03e-12 AS=3.69e-12 PD=1.934e-05 PS=9.82e-06
M73@2 N_CIN_M73@2_d N_U26_U36_drain_M73@2_g N_VDD_M73_s N_VDD_M79_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M73@3 N_CIN_M73@2_d N_U26_U36_drain_M73@3_g N_VDD_M73@3_s N_VDD_M79_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M73@4 N_CIN_M73@4_d N_U26_U36_drain_M73@4_g N_VDD_M73@3_s N_VDD_M79_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M79 N_U32_U1_nsgate_M79_d N_RENB_M79_g N_VDD_M79_s N_VDD_M79_b P18 L=2e-07
+ W=2.78e-06 AD=1.946e-12 AS=1.946e-12 PD=6.96e-06 PS=6.96e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M79_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M79_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M79_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M79_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D80 N_VSS_M19_b N_RENB_D80_neg DN18  AREA=1e-12 PJ=4e-06
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_VSSO_RM66_pos N_net_m66_VSSO_res_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
*
.include "pc3b25eu.dist.sp.PC3B25EU.pxi"
*
.ends
*
*
* File: pc3c01.dist.sp
* Created: Sun Jul  4 12:21:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c01.dist.sp.pex"
.subckt pc3c01  CCLK CP VDD VSS VDDO VSSO 
* 
M10 N_NODE_M10_d N_CCLK_M10_g N_VDD_M10_s N_VDD_M10_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M12 N_NODE_M10_d N_CCLK_M12_g N_VDD_M12_s N_VDD_M10_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M4 N_CP_M4_d N_NODE_M4_g N_VDD_M4_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M5 N_CP_M4_d N_NODE_M5_g N_VDD_M5_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M8 N_CP_M8_d N_NODE_M8_g N_VDD_M5_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M9 N_CP_M8_d N_NODE_M9_g N_VDD_M9_s N_VDD_M4_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D1 N_VSS_M11_b N_CCLK_D1_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M11 N_NODE_M11_d N_CCLK_M11_g N_VSS_M11_s N_VSS_M11_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M13 N_NODE_M11_d N_CCLK_M13_g N_VSS_M13_s N_VSS_M11_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M2 N_CP_M2_d N_NODE_M2_g N_VSS_M2_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M3 N_CP_M2_d N_NODE_M3_g N_VSS_M3_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_CP_M6_d N_NODE_M6_g N_VSS_M3_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M7 N_CP_M6_d N_NODE_M7_g N_VSS_M7_s N_VSS_M2_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
*
.include "pc3c01.dist.sp.PC3C01.pxi"
*
.ends
*
*
* File: pc3c02.dist.sp
* Created: Sun Jul  4 12:22:40 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c02.dist.sp.pex"
.subckt pc3c02  CCLK CP VDD VSS VDDO VSSO 
* 
M1 N_NODE_M1_d N_CCLK_M1_g N_VDD_M1_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_NODE_M1_d N_CCLK_M3_g N_VDD_M3_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M5 N_NODE_M5_d N_CCLK_M5_g N_VDD_M5_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M7 N_NODE_M5_d N_CCLK_M7_g N_VDD_M7_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M11 N_CP_M11_d N_NODE_M11_g N_VDD_M11_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M12 N_CP_M11_d N_NODE_M12_g N_VDD_M12_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M15 N_CP_M15_d N_NODE_M15_g N_VDD_M12_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M16 N_CP_M15_d N_NODE_M16_g N_VDD_M16_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M16_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M11_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D25 N_VSS_M2_b N_CCLK_D25_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M9 N_CP_M17_d N_NODE_M9_g N_VSS_M9_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M10 N_CP_M18_d N_NODE_M10_g N_VSS_M10_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M13 N_CP_M21_d N_NODE_M13_g N_VSS_M10_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_CP_M22_d N_NODE_M14_g N_VSS_M14_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M2 N_NODE_M2_d N_CCLK_M2_g N_VSS_M2_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4 N_NODE_M2_d N_CCLK_M4_g N_VSS_M4_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M17 N_CP_M17_d N_NODE_M17_g N_VSS_M17_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M18 N_CP_M18_d N_NODE_M18_g N_VSS_M17_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_NODE_M6_d N_CCLK_M6_g N_VSS_M6_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8 N_NODE_M6_d N_CCLK_M8_g N_VSS_M8_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M21 N_CP_M21_d N_NODE_M21_g N_VSS_M21_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M22_d N_NODE_M22_g N_VSS_M21_s N_VSS_M17_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c02.dist.sp.PC3C02.pxi"
*
.ends
*
*
* File: pc3c03.dist.sp
* Created: Sun Jul  4 12:22:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c03.dist.sp.pex"
.subckt pc3c03  CCLK CP VDD VSS VDDO VSSO 
* 
M17 N_CP_M33_d N_NODE_M17_g N_VSS_M17_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M18 N_CP_M34_d N_NODE_M18_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M21 N_CP_M37_d N_NODE_M21_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M38_d N_NODE_M22_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M25 N_CP_M41_d N_NODE_M25_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M26 N_CP_M42_d N_NODE_M26_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M29 N_CP_M45_d N_NODE_M29_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M30 N_CP_M46_d N_NODE_M30_g N_VSS_M30_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M1 N_NODE_M1_d N_CCLK_M1_g N_VDD_M1_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_NODE_M1_d N_CCLK_M3_g N_VDD_M3_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M5 N_NODE_M5_d N_CCLK_M5_g N_VDD_M5_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M7 N_NODE_M5_d N_CCLK_M7_g N_VDD_M7_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M9 N_NODE_M9_d N_CCLK_M9_g N_VDD_M9_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M11 N_NODE_M9_d N_CCLK_M11_g N_VDD_M11_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M13 N_NODE_M13_d N_CCLK_M13_g N_VDD_M13_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M15 N_NODE_M13_d N_CCLK_M15_g N_VDD_M15_s N_VDD_M1_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M19_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M27 N_CP_M27_d N_NODE_M27_g N_VDD_M24_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M28 N_CP_M27_d N_NODE_M28_g N_VDD_M28_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M31 N_CP_M31_d N_NODE_M31_g N_VDD_M28_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M32 N_CP_M31_d N_NODE_M32_g N_VDD_M32_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M35 N_CP_M35_d N_NODE_M35_g N_VDD_M32_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M36 N_CP_M35_d N_NODE_M36_g N_VDD_M36_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M39 N_CP_M39_d N_NODE_M39_g N_VDD_M36_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M40 N_CP_M39_d N_NODE_M40_g N_VDD_M40_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M43 N_CP_M43_d N_NODE_M43_g N_VDD_M40_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M44 N_CP_M43_d N_NODE_M44_g N_VDD_M44_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M47 N_CP_M47_d N_NODE_M47_g N_VDD_M44_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M48 N_CP_M47_d N_NODE_M48_g N_VDD_M48_s N_VDD_M19_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D49 N_VSS_M2_b N_CCLK_D49_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M2 N_NODE_M2_d N_CCLK_M2_g N_VSS_M2_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4 N_NODE_M2_d N_CCLK_M4_g N_VSS_M4_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M33 N_CP_M33_d N_NODE_M33_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M34 N_CP_M34_d N_NODE_M34_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_NODE_M6_d N_CCLK_M6_g N_VSS_M6_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M8 N_NODE_M6_d N_CCLK_M8_g N_VSS_M8_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_CP_M37_d N_NODE_M37_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M38 N_CP_M38_d N_NODE_M38_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M10 N_NODE_M10_d N_CCLK_M10_g N_VSS_M10_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M12 N_NODE_M10_d N_CCLK_M12_g N_VSS_M12_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41 N_CP_M41_d N_NODE_M41_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M42 N_CP_M42_d N_NODE_M42_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_NODE_M14_d N_CCLK_M14_g N_VSS_M14_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M16 N_NODE_M14_d N_CCLK_M16_g N_VSS_M16_s N_VSS_M2_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_CP_M45_d N_NODE_M45_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M46 N_CP_M46_d N_NODE_M46_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c03.dist.sp.PC3C03.pxi"
*
.ends
*
*
* File: pc3c04.dist.sp
* Created: Sun Jul  4 12:24:16 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3c04.dist.sp.pex"
.subckt pc3c04  CCLK CP VDD VSS VDDO VSSO 
* 
M1 N_CP_M33_d N_NODE_M1_g N_VSS_M1_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M2 N_CP_M34_d N_NODE_M2_g N_VSS_M2_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M5 N_CP_M37_d N_NODE_M5_g N_VSS_M2_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M6 N_CP_M38_d N_NODE_M6_g N_VSS_M6_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M9 N_CP_M41_d N_NODE_M9_g N_VSS_M6_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M10 N_CP_M42_d N_NODE_M10_g N_VSS_M10_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M13 N_CP_M45_d N_NODE_M13_g N_VSS_M10_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M14 N_CP_M46_d N_NODE_M14_g N_VSS_M14_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M17 N_CP_M49_d N_NODE_M17_g N_VSS_M14_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M18 N_CP_M50_d N_NODE_M18_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M21 N_CP_M53_d N_NODE_M21_g N_VSS_M18_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M22 N_CP_M54_d N_NODE_M22_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M25 N_CP_M57_d N_NODE_M25_g N_VSS_M22_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M26 N_CP_M58_d N_NODE_M26_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M29 N_CP_M61_d N_NODE_M29_g N_VSS_M26_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M30 N_CP_M62_d N_NODE_M30_g N_VSS_M30_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=9.869e-12 PD=1.49e-05 PS=2.922e-05
M65 N_NODE_M65_d N_CCLK_M65_g N_VDD_M65_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M67 N_NODE_M65_d N_CCLK_M67_g N_VDD_M67_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M69 N_NODE_M69_d N_CCLK_M69_g N_VDD_M69_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M71 N_NODE_M69_d N_CCLK_M71_g N_VDD_M71_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M73 N_NODE_M73_d N_CCLK_M73_g N_VDD_M73_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M75 N_NODE_M73_d N_CCLK_M75_g N_VDD_M75_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M77 N_NODE_M77_d N_CCLK_M77_g N_VDD_M77_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M79 N_NODE_M77_d N_CCLK_M79_g N_VDD_M79_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M81 N_NODE_M81_d N_CCLK_M81_g N_VDD_M81_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M83 N_NODE_M81_d N_CCLK_M83_g N_VDD_M83_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M85 N_NODE_M85_d N_CCLK_M85_g N_VDD_M85_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M87 N_NODE_M85_d N_CCLK_M87_g N_VDD_M87_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M89 N_NODE_M89_d N_CCLK_M89_g N_VDD_M89_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M91 N_NODE_M89_d N_CCLK_M91_g N_VDD_M91_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M93 N_NODE_M93_d N_CCLK_M93_g N_VDD_M93_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M95 N_NODE_M93_d N_CCLK_M95_g N_VDD_M95_s N_VDD_M65_b PHV L=3.6e-07 W=2.35e-05
+ AD=9.635e-12 AS=1.457e-11 PD=2.432e-05 PS=4.824e-05
M3 N_CP_M3_d N_NODE_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
M4 N_CP_M3_d N_NODE_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M7 N_CP_M7_d N_NODE_M7_g N_VDD_M4_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M8 N_CP_M7_d N_NODE_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M11 N_CP_M11_d N_NODE_M11_g N_VDD_M8_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M12 N_CP_M11_d N_NODE_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M15 N_CP_M15_d N_NODE_M15_g N_VDD_M12_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M16 N_CP_M15_d N_NODE_M16_g N_VDD_M16_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M19 N_CP_M19_d N_NODE_M19_g N_VDD_M16_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M20 N_CP_M19_d N_NODE_M20_g N_VDD_M20_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M23 N_CP_M23_d N_NODE_M23_g N_VDD_M20_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M24 N_CP_M23_d N_NODE_M24_g N_VDD_M24_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M27 N_CP_M27_d N_NODE_M27_g N_VDD_M24_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M28 N_CP_M27_d N_NODE_M28_g N_VDD_M28_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M31 N_CP_M31_d N_NODE_M31_g N_VDD_M28_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M32 N_CP_M31_d N_NODE_M32_g N_VDD_M32_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M35 N_CP_M35_d N_NODE_M35_g N_VDD_M32_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M36 N_CP_M35_d N_NODE_M36_g N_VDD_M36_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M39 N_CP_M39_d N_NODE_M39_g N_VDD_M36_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M40 N_CP_M39_d N_NODE_M40_g N_VDD_M40_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M43 N_CP_M43_d N_NODE_M43_g N_VDD_M40_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M44 N_CP_M43_d N_NODE_M44_g N_VDD_M44_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M47 N_CP_M47_d N_NODE_M47_g N_VDD_M44_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M48 N_CP_M47_d N_NODE_M48_g N_VDD_M48_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M51 N_CP_M51_d N_NODE_M51_g N_VDD_M48_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M52 N_CP_M51_d N_NODE_M52_g N_VDD_M52_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M55 N_CP_M55_d N_NODE_M55_g N_VDD_M52_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M56 N_CP_M55_d N_NODE_M56_g N_VDD_M56_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M59 N_CP_M59_d N_NODE_M59_g N_VDD_M56_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M60 N_CP_M59_d N_NODE_M60_g N_VDD_M60_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M63 N_CP_M63_d N_NODE_M63_g N_VDD_M60_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=1.617e-11 PD=3.334e-05 PS=3.334e-05
M64 N_CP_M63_d N_NODE_M64_g N_VDD_M64_s N_VDD_M3_b P18 L=1.8e-07 W=3.234e-05
+ AD=1.617e-11 AS=2.29614e-11 PD=3.334e-05 PS=6.61e-05
D97 N_VSS_M66_b N_CCLK_D97_neg DN18  AREA=4.624e-13 PJ=2.72e-06
M66 N_NODE_M66_d N_CCLK_M66_g N_VSS_M66_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M68 N_NODE_M66_d N_CCLK_M68_g N_VSS_M68_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M33 N_CP_M33_d N_NODE_M33_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M34 N_CP_M34_d N_NODE_M34_g N_VSS_M33_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M70 N_NODE_M70_d N_CCLK_M70_g N_VSS_M70_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M72 N_NODE_M70_d N_CCLK_M72_g N_VSS_M72_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_CP_M37_d N_NODE_M37_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M38 N_CP_M38_d N_NODE_M38_g N_VSS_M37_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M74 N_NODE_M74_d N_CCLK_M74_g N_VSS_M74_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M76 N_NODE_M74_d N_CCLK_M76_g N_VSS_M76_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41 N_CP_M41_d N_NODE_M41_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M42 N_CP_M42_d N_NODE_M42_g N_VSS_M41_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M78 N_NODE_M78_d N_CCLK_M78_g N_VSS_M78_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M80 N_NODE_M78_d N_CCLK_M80_g N_VSS_M80_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_CP_M45_d N_NODE_M45_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M46 N_CP_M46_d N_NODE_M46_g N_VSS_M45_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M82 N_NODE_M82_d N_CCLK_M82_g N_VSS_M82_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M84 N_NODE_M82_d N_CCLK_M84_g N_VSS_M84_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M49 N_CP_M49_d N_NODE_M49_g N_VSS_M49_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M50 N_CP_M50_d N_NODE_M50_g N_VSS_M49_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M86 N_NODE_M86_d N_CCLK_M86_g N_VSS_M86_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M88 N_NODE_M86_d N_CCLK_M88_g N_VSS_M88_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M53 N_CP_M53_d N_NODE_M53_g N_VSS_M53_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M54 N_CP_M54_d N_NODE_M54_g N_VSS_M53_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M90 N_NODE_M90_d N_CCLK_M90_g N_VSS_M90_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M92 N_NODE_M90_d N_CCLK_M92_g N_VSS_M92_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M57 N_CP_M57_d N_NODE_M57_g N_VSS_M57_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M58 N_CP_M58_d N_NODE_M58_g N_VSS_M57_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M94 N_NODE_M94_d N_CCLK_M94_g N_VSS_M94_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M96 N_NODE_M94_d N_CCLK_M96_g N_VSS_M96_s N_VSS_M66_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M61 N_CP_M61_d N_NODE_M61_g N_VSS_M61_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
M62 N_CP_M62_d N_NODE_M62_g N_VSS_M61_s N_VSS_M33_b N18 L=1.8e-07 W=1.39e-05
+ AD=6.95e-12 AS=6.95e-12 PD=1.49e-05 PS=1.49e-05
*
.include "pc3c04.dist.sp.PC3C04.pxi"
*
.ends
*
*
* File: pc3d00.dist.sp
* Created: Sun Jul  4 12:24:11 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d00.dist.sp.pex"
.subckt pc3d00  PAD PADR VDD VSS VDDO VSSO 
* 
M19 N_PAD_M25_d N_U18_U74$11_gate_M19_g N_VSSO_M19_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U18_U74$11_gate_M20_g N_VSSO_M20_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M21 N_PAD_M27_d N_U18_U74$11_gate_M21_g N_VSSO_M21_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M22 N_PAD_M28_d N_U18_U74$11_gate_M22_g N_VSSO_M19_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M29_d N_U18_U74$11_gate_M23_g N_VSSO_M23_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M24 N_PAD_M30_d N_U18_U74$11_gate_M24_g N_VSSO_M21_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
D32@2 N_VSS_D32@2_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@3 N_VSS_D32@3_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@4 N_VSS_D32@4_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@5 N_VSS_D32@5_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@6 N_VSS_D32@6_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32@7 N_VSS_D32@7_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D32 N_VSS_D32_pos N_VSSO_D32@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSSO_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSSO_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSSO_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSSO_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSSO_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSSO_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSSO_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XR15 N_VSS_R15_pos N_U18_U82_gate_R15_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR16 N_U18_U74$11_gate_R16_pos N_VSSO_R16_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR17 N_U18_U79$3_gate_R17_pos N_VDDO_R17_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M25 N_PAD_M25_d N_U18_U74$11_gate_M25_g N_VSSO_M25_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U18_U74$11_gate_M26_g N_VSSO_M25_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M27 N_PAD_M27_d N_U18_U74$11_gate_M27_g N_VSSO_M27_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M28 N_PAD_M28_d N_U18_U74$11_gate_M28_g N_VSSO_M27_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M29 N_PAD_M29_d N_U18_U74$11_gate_M29_g N_VSSO_M29_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M30 N_PAD_M30_d N_U18_U74$11_gate_M30_g N_VSSO_M29_s N_VSSO_M25_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR13 N_PADR_R13_pos N_noxref_2_R13_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR14 N_noxref_2_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M1 N_VDDO_M1_d N_U18_U79$3_gate_M1_g N_PAD_M1_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M2 N_VDDO_M5_d N_U18_U79$3_gate_M2_g N_PAD_M1_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_VDDO_M12_d N_U18_U79$3_gate_M3_g N_PAD_M3_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M4 N_VDDO_M4_d N_U18_U79$3_gate_M4_g N_PAD_M3_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M5 N_VDDO_M5_d N_U18_U79$3_gate_M5_g N_PAD_M5_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M6 N_VDDO_M6_d N_U18_U79$3_gate_M6_g N_PAD_M5_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M7 N_VDDO_M6_d N_U18_U79$3_gate_M7_g N_PAD_M7_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M8 N_VDDO_M8_d N_U18_U79$3_gate_M8_g N_PAD_M7_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M9 N_VDDO_M8_d N_U18_U79$3_gate_M9_g N_PAD_M9_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M10 N_VDDO_M10_d N_U18_U79$3_gate_M10_g N_PAD_M9_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M11 N_VDDO_M10_d N_U18_U79$3_gate_M11_g N_PAD_M11_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M12 N_VDDO_M12_d N_U18_U79$3_gate_M12_g N_PAD_M11_s N_VDDO_M5_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_PADR_M18_d N_U18_U82_gate_M18_g N_VSS_M18_s N_VSS_M18_b NHV L=4e-07
+ W=3e-05 AD=1.842e-10 AS=4.29e-11 PD=7.228e-05 PS=6.286e-05
*
.include "pc3d00.dist.sp.PC3D00.pxi"
*
.ends
*
*
* File: pc3d01d.dist.sp
* Created: Sun Jul  4 12:26:04 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d01d.dist.sp.pex"
.subckt pc3d01d  CIN PAD VDD VSS VDDO VSSO 
* 
M1 N_U14_padr_M1_d N_net_m1_VDDO_res_M1_g U15_U22_source N_VSS_M12_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M2 U15_U22_source N_net_m2_VDDO_res_M2_g N_VSSO_M2_s N_VSS_M12_b NHV L=5.5e-06
+ W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M16 N_PAD_M22_d N_U14_MN4$11_gate_M16_g N_VSSO_M16_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M23_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M18 N_PAD_M24_d N_U14_MN4$11_gate_M18_g N_VSSO_M18_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M25_d N_U14_MN4$11_gate_M19_g N_VSSO_M16_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U14_MN4$11_gate_M20_g N_VSSO_M20_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M21 N_PAD_M27_d N_U14_MN4$11_gate_M21_g N_VSSO_M18_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR28 N_U14_MN4$11_gate_R28_pos N_VSSO_R28_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VDDO_res_RM1_pos N_VDDO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_VDDO_RM1_neg N_net_m2_VDDO_res_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
M22 N_PAD_M22_d N_U14_MN4$11_gate_M22_g N_VSSO_M22_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M23 N_PAD_M23_d N_U14_MN4$11_gate_M23_g N_VSSO_M22_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U14_MN4$11_gate_M24_g N_VSSO_M24_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U14_MN4$11_gate_M25_g N_VSSO_M24_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U14_MN4$11_gate_M26_g N_VSSO_M26_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M27 N_PAD_M27_d N_U14_MN4$11_gate_M27_g N_VSSO_M26_s N_VSSO_M22_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M30 N_VDDO_M33_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M40_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M33 N_VDDO_M33_d N_U14_pgate_tol_M33_g N_PAD_M33_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U14_pgate_tol_M34_g N_PAD_M33_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_VDDO_M34_d N_U14_pgate_tol_M35_g N_PAD_M35_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U14_pgate_tol_M36_g N_PAD_M35_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_VDDO_M36_d N_U14_pgate_tol_M37_g N_PAD_M37_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_VDDO_M38_d N_U14_pgate_tol_M38_g N_PAD_M37_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M39 N_VDDO_M38_d N_U14_pgate_tol_M39_g N_PAD_M39_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M40 N_VDDO_M40_d N_U14_pgate_tol_M40_g N_PAD_M39_s N_VDDO_M33_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR14 N_X28/noxref_9_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR15 N_X28/noxref_9_R15_pos N_U14_padr_R15_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M12 N_U14_pgate_tol_M12_s N_net_m12_VDDO_res_M12_g N_U14_pgate_tol_M12_s
+ N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M12@2 N_U14_pgate_tol_M12@2_s N_net_m12_VDDO_res_M12@2_g
+ N_U14_pgate_tol_M12@2_s N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M12@3 N_U14_pgate_tol_M12@3_s N_net_m12_VDDO_res_M12@3_g
+ N_U14_pgate_tol_M12@3_s N_VSS_M12_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M10 N_VDDO_M10_d N_net_m10_VDDO_res_M10_g N_U14_pgate_tol_M10_s N_VSS_M12_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M8 N_U14_padr_M8_d N_net_m8_VSSO_res_M8_g N_VSSO_M8_s N_VSS_M12_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_U14_padr_M8@2_d N_net_m8_VSSO_res_M8@2_g N_VSSO_M8_s N_VSS_M12_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7 N_U9_MPI1_drain_M7_d N_U14_padr_M7_g N_VSSO_M7_s N_VSS_M12_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M9 N_CIN_M9_d N_U9_MPI1_drain_M9_g N_VSS_M9_s N_VSS_M12_b NHV L=3.6e-07 W=6e-06
+ AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M13 N_U14_pgate_tol_M13_s N_net_m13_VSSO_res_M13_g N_U14_pgate_tol_M13_s
+ N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11
+ PD=1.749e-05 PS=3.458e-05
M13@2 N_U14_pgate_tol_M13@2_s N_net_m13_VSSO_res_M13@2_g
+ N_U14_pgate_tol_M13@2_s N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12
+ AS=6.8347e-12 PD=1.749e-05 PS=1.749e-05
M13@3 N_U14_pgate_tol_M13@3_s N_net_m13_VSSO_res_M13@3_g
+ N_U14_pgate_tol_M13@3_s N_VDDO_M13_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11
+ AS=6.8347e-12 PD=3.46e-05 PS=1.749e-05
M11 N_U14_pgate_tol_M11_d N_net_m11_VSSO_res_M11_g N_VDDO_M11_s N_VDDO_M13_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M5 N_U14_padr_M5_d N_net_m5_VDDO_res_M5_g N_VDDO_M5_s N_VDDO_M13_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 U9_MPI2_drain N_U14_padr_M3_g N_VDDO_M3_s N_VDDO_M13_b PHV L=3.6e-07 W=2e-05
+ AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M4 N_U9_MPI1_drain_M4_d N_U14_padr_M4_g U9_MPI2_drain N_VDDO_M13_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M6 N_CIN_M6_d N_U9_MPI1_drain_M6_g N_VDD_M6_s N_VDD_M6_b PHV L=3.6e-07 W=8e-06
+ AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M6@2 N_CIN_M6@2_d N_U9_MPI1_drain_M6@2_g N_VDD_M6_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M6@3 N_CIN_M6@2_d N_U9_MPI1_drain_M6@3_g N_VDD_M6@3_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M6@4 N_CIN_M6@4_d N_U9_MPI1_drain_M6@4_g N_VDD_M6@3_s N_VDD_M6_b PHV L=3.6e-07
+ W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM5 N_net_m5_VDDO_res_RM5_pos N_VDDO_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM13 N_VSSO_RM13_pos N_net_m13_VSSO_res_RM13_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM12 N_VDDO_RM12_pos N_net_m12_VDDO_res_RM12_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM10 N_VDDO_RM10_pos N_net_m10_VDDO_res_RM10_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM11 N_net_m11_VSSO_res_RM11_pos N_VSSO_RM11_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM8 N_VSSO_RM8_pos N_net_m8_VSSO_res_RM8_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U9_MPI2_drain 0 0.0173376f
*
.include "pc3d01d.dist.sp.PC3D01D.pxi"
*
.ends
*
*
* File: pc3d01.dist.sp
* Created: Sun Jul  4 12:26:00 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d01.dist.sp.pex"
.subckt pc3d01  CIN PAD VDD VSS VDDO VSSO 
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X24/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X24/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M37 N_U14_padr_M37_d N_net_m37_VSSO_res_M37_g N_VSSO_M37_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M37@2 N_U14_padr_M37@2_d N_net_m37_VSSO_res_M37@2_g N_VSSO_M37_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36 N_U9_MPI1_drain_M36_d N_U14_padr_M36_g N_VSSO_M36_s N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M38 N_CIN_M38_d N_U9_MPI1_drain_M38_g N_VSS_M38_s N_VSS_M3_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M34 N_U14_padr_M34_d N_net_m34_VDDO_res_M34_g N_VDDO_M34_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M32 U9_MPI2_drain N_U14_padr_M32_g N_VDDO_M32_s N_VDDO_M4_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M33 N_U9_MPI1_drain_M33_d N_U14_padr_M33_g U9_MPI2_drain N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M35 N_CIN_M35_d N_U9_MPI1_drain_M35_g N_VDD_M35_s N_VDD_M35_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M35@2 N_CIN_M35@2_d N_U9_MPI1_drain_M35@2_g N_VDD_M35_s N_VDD_M35_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M35@3 N_CIN_M35@2_d N_U9_MPI1_drain_M35@3_g N_VDD_M35@3_s N_VDD_M35_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M35@4 N_CIN_M35@4_d N_U9_MPI1_drain_M35@4_g N_VDD_M35@3_s N_VDD_M35_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM34 N_net_m34_VDDO_res_RM34_pos N_VDDO_RM34_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U9_MPI2_drain 0 0.0173376f
*
.include "pc3d01.dist.sp.PC3D01.pxi"
*
.ends
*
*
* File: pc3d01u.dist.sp
* Created: Sun Jul  4 12:27:46 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d01u.dist.sp.pex"
.subckt pc3d01u  CIN PAD VDD VSS VDDO VSSO 
* 
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M12_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M19_d N_U14_MN4$11_gate_M13_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U14_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M5_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR20 N_U14_MN4$11_gate_R20_pos N_VSSO_R20_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M19_d N_U14_MN4$11_gate_M19_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
M21 N_VDDO_M21_d N_U14_pgate_tol_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M22 N_VDDO_M25_d N_U14_pgate_tol_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_U14_pgate_tol_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U14_pgate_tol_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U14_pgate_tol_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U14_pgate_tol_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR6 N_X26/noxref_9_R6_pos N_PAD_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR7 N_X26/noxref_9_R7_pos N_U14_padr_R7_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M4 N_U14_pgate_tol_M4_s N_net_m4_VDDO_res_M4_g N_U14_pgate_tol_M4_s N_VSS_M4_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VDDO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VDDO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_VDDO_M2_d N_net_m2_VDDO_res_M2_g N_U14_pgate_tol_M2_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U14_padr_M38_d N_net_m38_VSSO_res_M38_g N_VSSO_M38_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U14_padr_M38@2_d N_net_m38_VSSO_res_M38@2_g N_VSSO_M38_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M37 N_U9_MPI1_drain_M37_d N_U14_padr_M37_g N_VSSO_M37_s N_VSS_M4_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M39 N_CIN_M39_d N_U9_MPI1_drain_M39_g N_VSS_M39_s N_VSS_M4_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M5 N_U14_pgate_tol_M5_s N_net_m5_VSSO_res_M5_g N_U14_pgate_tol_M5_s N_VDDO_M5_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M5@2 N_U14_pgate_tol_M5@2_s N_net_m5_VSSO_res_M5@2_g N_U14_pgate_tol_M5@2_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M5@3 N_U14_pgate_tol_M5@3_s N_net_m5_VSSO_res_M5@3_g N_U14_pgate_tol_M5@3_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M3 N_U14_pgate_tol_M3_d N_net_m3_VSSO_res_M3_g N_VDDO_M3_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M35 N_U14_padr_M35_d N_net_m35_VDDO_res_M35_g N_VDDO_M35_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M33 U9_MPI2_drain N_U14_padr_M33_g N_VDDO_M33_s N_VDDO_M5_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M34 N_U9_MPI1_drain_M34_d N_U14_padr_M34_g U9_MPI2_drain N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M36 N_CIN_M36_d N_U9_MPI1_drain_M36_g N_VDD_M36_s N_VDD_M36_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M36@2 N_CIN_M36@2_d N_U9_MPI1_drain_M36@2_g N_VDD_M36_s N_VDD_M36_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M36@3 N_CIN_M36@2_d N_U9_MPI1_drain_M36@3_g N_VDD_M36@3_s N_VDD_M36_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M36@4 N_CIN_M36@4_d N_U9_MPI1_drain_M36@4_g N_VDD_M36@3_s N_VDD_M36_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM35 N_net_m35_VDDO_res_RM35_pos N_VDDO_RM35_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM5 N_VSSO_RM5_pos N_net_m5_VSSO_res_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM4 N_VDDO_RM4_pos N_net_m4_VDDO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_VDDO_RM2_pos N_net_m2_VDDO_res_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_net_m3_VSSO_res_RM3_pos N_VSSO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM38 N_VSSO_RM38_pos N_net_m38_VSSO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U9_MPI2_drain 0 0.0173376f
*
.include "pc3d01u.dist.sp.PC3D01U.pxi"
*
.ends
*
*
* File: pc3d11d.dist.sp
* Created: Sun Jul  4 12:29:18 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d11d.dist.sp.pex"
.subckt pc3d11d  CIN PAD VDD VSS VDDO VSSO 
* 
M32 N_U14_padr_M32_d N_net_m32_VDDO_res_M32_g U15_U22_source N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M33 U15_U22_source N_net_m33_VDDO_res_M33_g N_VSSO_M33_s N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM32 N_net_m32_VDDO_res_RM32_pos N_VDDO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM33 N_VDDO_RM32_neg N_net_m33_VDDO_res_RM33_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X28/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X28/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_U14_padr_M39_d N_net_m39_VSSO_res_M39_g N_VSSO_M39_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U14_padr_M39@2_d N_net_m39_VSSO_res_M39@2_g N_VSSO_M39_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40 N_U9_MNI1_drain_M40_d N_U14_padr_M40_g N_VSSO_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M41 N_CIN_M41_d N_U9_U19_gate_M41_g N_VSS_M41_s N_VSS_M3_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M42 N_U9_U19_gate_M42_d N_U9_MNI1_drain_M42_g N_VSSO_M42_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1.5e-05 AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M34 N_U14_padr_M34_d N_net_m34_VDDO_res_M34_g N_VDDO_M34_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M36 U9_MPI1_source N_U14_padr_M36_g N_VDDO_M36_s N_VDDO_M4_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M35 N_U9_MNI1_drain_M35_d N_U14_padr_M35_g U9_MPI1_source N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M37 N_U9_U19_gate_M37_d N_U9_MNI1_drain_M37_g N_VDDO_M37_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M37@2 N_U9_U19_gate_M37_d N_U9_MNI1_drain_M37@2_g N_VDDO_M37@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M38 N_CIN_M38_d N_U9_U19_gate_M38_g N_VDD_M38_s N_VDD_M38_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M38@2 N_CIN_M38@2_d N_U9_U19_gate_M38@2_g N_VDD_M38_s N_VDD_M38_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M38@3 N_CIN_M38@2_d N_U9_U19_gate_M38@3_g N_VDD_M38@3_s N_VDD_M38_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M38@4 N_CIN_M38@4_d N_U9_U19_gate_M38@4_g N_VDD_M38@3_s N_VDD_M38_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM34 N_net_m34_VDDO_res_RM34_pos N_VDDO_RM34_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U9_MPI1_source 0 0.0173376f
*
.include "pc3d11d.dist.sp.PC3D11D.pxi"
*
.ends
*
*
* File: pc3d11.dist.sp
* Created: Sun Jul  4 12:27:41 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d11.dist.sp.pex"
.subckt pc3d11  CIN PAD VDD VSS VDDO VSSO 
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X24/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X24/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M37 N_U14_padr_M37_d N_net_m37_VSSO_res_M37_g N_VSSO_M37_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M37@2 N_U14_padr_M37@2_d N_net_m37_VSSO_res_M37@2_g N_VSSO_M37_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38 N_U9_MNI1_drain_M38_d N_U14_padr_M38_g N_VSSO_M38_s N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M39 N_CIN_M39_d N_U9_U19_gate_M39_g N_VSS_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M40 N_U9_U19_gate_M40_d N_U9_MNI1_drain_M40_g N_VSSO_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1.5e-05 AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M32 N_U14_padr_M32_d N_net_m32_VDDO_res_M32_g N_VDDO_M32_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M34 U9_MPI1_source N_U14_padr_M34_g N_VDDO_M34_s N_VDDO_M4_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M33 N_U9_MNI1_drain_M33_d N_U14_padr_M33_g U9_MPI1_source N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M35 N_U9_U19_gate_M35_d N_U9_MNI1_drain_M35_g N_VDDO_M35_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M35@2 N_U9_U19_gate_M35_d N_U9_MNI1_drain_M35@2_g N_VDDO_M35@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M36 N_CIN_M36_d N_U9_U19_gate_M36_g N_VDD_M36_s N_VDD_M36_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M36@2 N_CIN_M36@2_d N_U9_U19_gate_M36@2_g N_VDD_M36_s N_VDD_M36_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M36@3 N_CIN_M36@2_d N_U9_U19_gate_M36@3_g N_VDD_M36@3_s N_VDD_M36_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M36@4 N_CIN_M36@4_d N_U9_U19_gate_M36@4_g N_VDD_M36@3_s N_VDD_M36_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM32 N_net_m32_VDDO_res_RM32_pos N_VDDO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U9_MPI1_source 0 0.0173376f
*
.include "pc3d11.dist.sp.PC3D11.pxi"
*
.ends
*
*
* File: pc3d11u.dist.sp
* Created: Sun Jul  4 12:29:17 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d11u.dist.sp.pex"
.subckt pc3d11u  CIN PAD VDD VSS VDDO VSSO 
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U14_padr_M32_d N_net_m32_VSSO_res_M32_g N_VDDO_M32_s N_VDDO_M4_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X26/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X26/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U14_padr_M38_d N_net_m38_VSSO_res_M38_g N_VSSO_M38_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U14_padr_M38@2_d N_net_m38_VSSO_res_M38@2_g N_VSSO_M38_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U9_MNI1_drain_M39_d N_U14_padr_M39_g N_VSSO_M39_s N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M40 N_CIN_M40_d N_U9_U19_gate_M40_g N_VSS_M40_s N_VSS_M3_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M41 N_U9_U19_gate_M41_d N_U9_MNI1_drain_M41_g N_VSSO_M41_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1.5e-05 AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M33 N_U14_padr_M33_d N_net_m33_VDDO_res_M33_g N_VDDO_M33_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M35 U9_MPI1_source N_U14_padr_M35_g N_VDDO_M35_s N_VDDO_M4_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M34 N_U9_MNI1_drain_M34_d N_U14_padr_M34_g U9_MPI1_source N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M36 N_U9_U19_gate_M36_d N_U9_MNI1_drain_M36_g N_VDDO_M36_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M36@2 N_U9_U19_gate_M36_d N_U9_MNI1_drain_M36@2_g N_VDDO_M36@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M37 N_CIN_M37_d N_U9_U19_gate_M37_g N_VDD_M37_s N_VDD_M37_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M37@2 N_CIN_M37@2_d N_U9_U19_gate_M37@2_g N_VDD_M37_s N_VDD_M37_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M37@3 N_CIN_M37@2_d N_U9_U19_gate_M37@3_g N_VDD_M37@3_s N_VDD_M37_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M37@4 N_CIN_M37@4_d N_U9_U19_gate_M37@4_g N_VDD_M37@3_s N_VDD_M37_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
XRM33 N_net_m33_VDDO_res_RM33_pos N_VDDO_RM33_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM38 N_VSSO_RM38_pos N_net_m38_VSSO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U9_MPI1_source 0 0.0173376f
*
.include "pc3d11u.dist.sp.PC3D11U.pxi"
*
.ends
*
*
* File: pc3d21d.dist.sp
* Created: Sun Jul  4 12:30:51 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d21d.dist.sp.pex"
.subckt pc3d21d  CIN PAD VDD VSS VDDO VSSO 
* 
M32 N_U14_padr_M32_d N_net_m32_VDDO_res_M32_g U15_U22_source N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M33 U15_U22_source N_net_m33_VDDO_res_M33_g N_VSSO_M33_s N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM32 N_net_m32_VDDO_res_RM32_pos N_VDDO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM33 N_VDDO_RM32_neg N_net_m33_VDDO_res_RM33_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X28/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X28/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U14_padr_M36_d N_net_m36_VSSO_res_M36_g N_VSSO_M36_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36@2 N_U14_padr_M36@2_d N_net_m36_VSSO_res_M36@2_g N_VSSO_M36_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M34 N_U9_U34_drain_M34_d N_U14_padr_M34_g N_VSSO_M34_s N_VSS_M3_b NHV L=3.6e-07
+ W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M35 N_U9_U36_drain_M35_d N_U14_padr_M35_g N_U9_U34_drain_M34_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M37 N_VDDO_M37_d N_U9_U36_drain_M37_g N_U9_U34_drain_M37_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M38 N_CIN_M38_d N_U9_U36_drain_M38_g N_VSS_M38_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M41 N_U14_padr_M41_d N_net_m41_VDDO_res_M41_g N_VDDO_M41_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U14_padr_M41_d N_net_m41_VDDO_res_M41@2_g N_VDDO_M41@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40 N_U9_U30_source_M40_d N_U14_padr_M40_g N_VDDO_M40_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M39 N_U9_U36_drain_M39_d N_U14_padr_M39_g N_U9_U30_source_M40_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M42 N_VSSO_M42_d N_U9_U36_drain_M42_g N_U9_U30_source_M42_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M43 N_CIN_M43_d N_U9_U36_drain_M43_g N_VDD_M43_s N_VDD_M43_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M43@2 N_CIN_M43@2_d N_U9_U36_drain_M43@2_g N_VDD_M43_s N_VDD_M43_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M43@3 N_CIN_M43@2_d N_U9_U36_drain_M43@3_g N_VDD_M43@3_s N_VDD_M43_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M43@4 N_CIN_M43@4_d N_U9_U36_drain_M43@4_g N_VDD_M43@3_s N_VDD_M43_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM41 N_net_m41_VDDO_res_RM41_pos N_VDDO_RM41_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM36 N_VSSO_RM36_pos N_net_m36_VSSO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d21d.dist.sp.PC3D21D.pxi"
*
.ends
*
*
* File: pc3d21eu.dist.sp
* Created: Sun Jul  4 12:32:30 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d21eu.dist.sp.pex"
.subckt pc3d21eu  CIN PAD RENB VDD VSS VDDO VSSO 
* 
M46 N_U17_U1_OUTSHIFT_M46_d N_U17_U1_nsgate_M46_g N_VSSO_M46_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M45 N_U17_U1_U6_drain_M45_d N_RENB_M45_g N_VSSO_M45_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_U17_U1_nsgate_M42_d N_RENB_M42_g N_VSS_M42_s N_VSS_M3_b N18 L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M49 N_U14_padr_M49_d N_U17_U1_OUTSHIFT_M49_g N_VDDO_M49_s N_VDDO_M4_b PHV
+ L=2e-06 W=2e-06 AD=4.26e-12 AS=4.24e-12 PD=8.26e-06 PS=8.24e-06
M43 N_U17_U1_U6_drain_M43_d N_U17_U1_OUTSHIFT_M43_g N_VDDO_M43_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
M44 N_U17_U1_OUTSHIFT_M44_d N_U17_U1_U6_drain_M44_g N_VDDO_M43_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=6e-06 AD=3.72e-12 AS=2.46e-12 PD=1.324e-05 PS=6.82e-06
M47 N_U17_U1_nsgate_M47_d N_RENB_M47_g N_VDD_M47_s N_VDD_M41_b P18 L=2e-07
+ W=2.78e-06 AD=1.946e-12 AS=1.946e-12 PD=6.96e-06 PS=6.96e-06
D48 N_VSS_M3_b N_RENB_D48_neg DN18  AREA=1e-12 PJ=4e-06
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X32/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X32/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U14_padr_M34_d N_net_m34_VSSO_res_M34_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M34@2 N_U14_padr_M34@2_d N_net_m34_VSSO_res_M34@2_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M32 N_U9_U34_drain_M32_d N_U14_padr_M32_g N_VSSO_M32_s N_VSS_M3_b NHV L=3.6e-07
+ W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M33 N_U9_U36_drain_M33_d N_U14_padr_M33_g N_U9_U34_drain_M32_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M35 N_VDDO_M35_d N_U9_U36_drain_M35_g N_U9_U34_drain_M35_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M36 N_CIN_M36_d N_U9_U36_drain_M36_g N_VSS_M36_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M39 N_U14_padr_M39_d N_net_m39_VDDO_res_M39_g N_VDDO_M39_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M38 N_U9_U30_source_M38_d N_U14_padr_M38_g N_VDDO_M38_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M37 N_U9_U36_drain_M37_d N_U14_padr_M37_g N_U9_U30_source_M38_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M40 N_VSSO_M40_d N_U9_U36_drain_M40_g N_U9_U30_source_M40_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M41 N_CIN_M41_d N_U9_U36_drain_M41_g N_VDD_M41_s N_VDD_M41_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M41@2 N_CIN_M41@2_d N_U9_U36_drain_M41@2_g N_VDD_M41_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@3 N_CIN_M41@2_d N_U9_U36_drain_M41@3_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@4 N_CIN_M41@4_d N_U9_U36_drain_M41@4_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM39 N_net_m39_VDDO_res_RM39_pos N_VDDO_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM34 N_VSSO_RM34_pos N_net_m34_VSSO_res_RM34_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d21eu.dist.sp.PC3D21EU.pxi"
*
.ends
*
*
* File: pc3d21.dist.sp
* Created: Sun Jul  4 12:31:01 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d21.dist.sp.pex"
.subckt pc3d21  CIN PAD VDD VSS VDDO VSSO 
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X24/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X24/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U14_padr_M34_d N_net_m34_VSSO_res_M34_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M34@2 N_U14_padr_M34@2_d N_net_m34_VSSO_res_M34@2_g N_VSSO_M34_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M32 N_U9_U34_drain_M32_d N_U14_padr_M32_g N_VSSO_M32_s N_VSS_M3_b NHV L=3.6e-07
+ W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M33 N_U9_U36_drain_M33_d N_U14_padr_M33_g N_U9_U34_drain_M32_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M35 N_VDDO_M35_d N_U9_U36_drain_M35_g N_U9_U34_drain_M35_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M36 N_CIN_M36_d N_U9_U36_drain_M36_g N_VSS_M36_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M39 N_U14_padr_M39_d N_net_m39_VDDO_res_M39_g N_VDDO_M39_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M39@2 N_U14_padr_M39_d N_net_m39_VDDO_res_M39@2_g N_VDDO_M39@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38 N_U9_U30_source_M38_d N_U14_padr_M38_g N_VDDO_M38_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M37 N_U9_U36_drain_M37_d N_U14_padr_M37_g N_U9_U30_source_M38_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M40 N_VSSO_M40_d N_U9_U36_drain_M40_g N_U9_U30_source_M40_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M41 N_CIN_M41_d N_U9_U36_drain_M41_g N_VDD_M41_s N_VDD_M41_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M41@2 N_CIN_M41@2_d N_U9_U36_drain_M41@2_g N_VDD_M41_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@3 N_CIN_M41@2_d N_U9_U36_drain_M41@3_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M41@4 N_CIN_M41@4_d N_U9_U36_drain_M41@4_g N_VDD_M41@3_s N_VDD_M41_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM39 N_net_m39_VDDO_res_RM39_pos N_VDDO_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM34 N_VSSO_RM34_pos N_net_m34_VSSO_res_RM34_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d21.dist.sp.PC3D21.pxi"
*
.ends
*
*
* File: pc3d21u.dist.sp
* Created: Sun Jul  4 12:32:31 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d21u.dist.sp.pex"
.subckt pc3d21u  CIN PAD VDD VSS VDDO VSSO 
* 
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M12_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M19_d N_U14_MN4$11_gate_M13_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U14_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M5_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR20 N_U14_MN4$11_gate_R20_pos N_VSSO_R20_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M19_d N_U14_MN4$11_gate_M19_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
M21 N_VDDO_M21_d N_U14_pgate_tol_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M22 N_VDDO_M25_d N_U14_pgate_tol_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_U14_pgate_tol_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U14_pgate_tol_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U14_pgate_tol_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U14_pgate_tol_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR6 N_X26/noxref_9_R6_pos N_PAD_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR7 N_X26/noxref_9_R7_pos N_U14_padr_R7_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M4 N_U14_pgate_tol_M4_s N_net_m4_VDDO_res_M4_g N_U14_pgate_tol_M4_s N_VSS_M4_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VDDO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VDDO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_VDDO_M2_d N_net_m2_VDDO_res_M2_g N_U14_pgate_tol_M2_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M35 N_U14_padr_M35_d N_net_m35_VSSO_res_M35_g N_VSSO_M35_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M35@2 N_U14_padr_M35@2_d N_net_m35_VSSO_res_M35@2_g N_VSSO_M35_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33 N_U9_U34_drain_M33_d N_U14_padr_M33_g N_VSSO_M33_s N_VSS_M4_b NHV L=3.6e-07
+ W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M34 N_U9_U36_drain_M34_d N_U14_padr_M34_g N_U9_U34_drain_M33_d N_VSS_M4_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M36 N_VDDO_M36_d N_U9_U36_drain_M36_g N_U9_U34_drain_M36_s N_VSS_M4_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M37 N_CIN_M37_d N_U9_U36_drain_M37_g N_VSS_M37_s N_VSS_M4_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M5 N_U14_pgate_tol_M5_s N_net_m5_VSSO_res_M5_g N_U14_pgate_tol_M5_s N_VDDO_M5_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M5@2 N_U14_pgate_tol_M5@2_s N_net_m5_VSSO_res_M5@2_g N_U14_pgate_tol_M5@2_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M5@3 N_U14_pgate_tol_M5@3_s N_net_m5_VSSO_res_M5@3_g N_U14_pgate_tol_M5@3_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M3 N_U14_pgate_tol_M3_d N_net_m3_VSSO_res_M3_g N_VDDO_M3_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M40 N_U14_padr_M40_d N_net_m40_VDDO_res_M40_g N_VDDO_M40_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U14_padr_M40_d N_net_m40_VDDO_res_M40@2_g N_VDDO_M40@2_s N_VDDO_M5_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M39 N_U9_U30_source_M39_d N_U14_padr_M39_g N_VDDO_M39_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M38 N_U9_U36_drain_M38_d N_U14_padr_M38_g N_U9_U30_source_M39_d N_VDDO_M5_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M41 N_VSSO_M41_d N_U9_U36_drain_M41_g N_U9_U30_source_M41_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M42 N_CIN_M42_d N_U9_U36_drain_M42_g N_VDD_M42_s N_VDD_M42_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M42@2 N_CIN_M42@2_d N_U9_U36_drain_M42@2_g N_VDD_M42_s N_VDD_M42_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M42@3 N_CIN_M42@2_d N_U9_U36_drain_M42@3_g N_VDD_M42@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M42@4 N_CIN_M42@4_d N_U9_U36_drain_M42@4_g N_VDD_M42@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM5 N_VSSO_RM5_pos N_net_m5_VSSO_res_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM4 N_VDDO_RM4_pos N_net_m4_VDDO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_VDDO_RM2_pos N_net_m2_VDDO_res_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_net_m3_VSSO_res_RM3_pos N_VSSO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM35 N_VSSO_RM35_pos N_net_m35_VSSO_res_RM35_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d21u.dist.sp.PC3D21U.pxi"
*
.ends
*
*
* File: pc3d31d.dist.sp
* Created: Sun Jul  4 12:34:21 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d31d.dist.sp.pex"
.subckt pc3d31d  CIN PAD VDD VSS VDDO VSSO 
* 
M32 N_U14_padr_M32_d N_net_m32_VDDO_res_M32_g U15_U22_source N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M33 U15_U22_source N_net_m33_VDDO_res_M33_g N_VSSO_M33_s N_VSS_M3_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM32 N_net_m32_VDDO_res_RM32_pos N_VDDO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM33 N_VDDO_RM32_neg N_net_m33_VDDO_res_RM33_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X28/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X28/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M43 N_U14_padr_M43_d N_net_m43_VSSO_res_M43_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U14_padr_M43@2_d N_net_m43_VSSO_res_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U9_U33_source_M41_d N_U14_padr_M41_g N_VSSO_M41_s N_VSS_M3_b NHV
+ L=3.6e-07 W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M42 N_U9_U41_gate_M42_d N_U14_padr_M42_g N_U9_U33_source_M41_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M40 N_VDDO_M40_d N_U9_U41_gate_M40_g N_U9_U33_source_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M44 N_U9_U43_drain_M44_d N_U9_U41_gate_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M44@2 N_U9_U43_drain_M44_d N_U9_U41_gate_M44@2_g N_VSSO_M44@2_s N_VSS_M3_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M45 N_CIN_M45_d N_U9_U43_drain_M45_g N_VSS_M45_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M37 N_U14_padr_M37_d N_net_m37_VDDO_res_M37_g N_VDDO_M37_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37@2 N_U14_padr_M37_d N_net_m37_VDDO_res_M37@2_g N_VDDO_M37@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M36 N_U9_U41_source_M36_d N_U14_padr_M36_g N_VDDO_M36_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M35 N_U9_U41_gate_M35_d N_U14_padr_M35_g N_U9_U41_source_M36_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M34 N_VSSO_M34_d N_U9_U41_gate_M34_g N_U9_U41_source_M34_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M38 N_U9_U43_drain_M38_d N_U9_U41_gate_M38_g N_VDDO_M38_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M38@2 N_U9_U43_drain_M38_d N_U9_U41_gate_M38@2_g N_VDDO_M38@2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M39 N_CIN_M39_d N_U9_U43_drain_M39_g N_VDD_M39_s N_VDD_M39_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M39@2 N_CIN_M39@2_d N_U9_U43_drain_M39@2_g N_VDD_M39_s N_VDD_M39_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M39@3 N_CIN_M39@2_d N_U9_U43_drain_M39@3_g N_VDD_M39@3_s N_VDD_M39_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M39@4 N_CIN_M39@4_d N_U9_U43_drain_M39@4_g N_VDD_M39@3_s N_VDD_M39_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM37 N_net_m37_VDDO_res_RM37_pos N_VDDO_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM43 N_VSSO_RM43_pos N_net_m43_VSSO_res_RM43_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d31d.dist.sp.PC3D31D.pxi"
*
.ends
*
*
* File: pc3d31.dist.sp
* Created: Sun Jul  4 12:34:24 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d31.dist.sp.pex"
.subckt pc3d31  CIN PAD VDD VSS VDDO VSSO 
* 
M7 N_PAD_M13_d N_U14_MN4$11_gate_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M11_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 N_U14_MN4$11_gate_R19_pos N_VSSO_R19_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M13 N_PAD_M13_d N_U14_MN4$11_gate_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M17_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_VDDO_M20_d N_U14_pgate_tol_M20_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M21 N_VDDO_M24_d N_U14_pgate_tol_M21_g N_PAD_M20_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M31_d N_U14_pgate_tol_M22_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M23_d N_U14_pgate_tol_M23_g N_PAD_M22_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M24_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M25_d N_U14_pgate_tol_M26_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M27_d N_U14_pgate_tol_M27_g N_PAD_M26_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M27_d N_U14_pgate_tol_M28_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M29_d N_U14_pgate_tol_M29_g N_PAD_M28_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M29_d N_U14_pgate_tol_M30_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M31_d N_U14_pgate_tol_M31_g N_PAD_M30_s N_VDDO_M24_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR5 N_X24/noxref_9_R5_pos N_PAD_R5_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR6 N_X24/noxref_9_R6_pos N_U14_padr_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M3 N_U14_pgate_tol_M3_s N_net_m3_VDDO_res_M3_g N_U14_pgate_tol_M3_s N_VSS_M3_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M3@2 N_U14_pgate_tol_M3@2_s N_net_m3_VDDO_res_M3@2_g N_U14_pgate_tol_M3@2_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M3@3 N_U14_pgate_tol_M3@3_s N_net_m3_VDDO_res_M3@3_g N_U14_pgate_tol_M3@3_s
+ N_VSS_M3_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M1 N_VDDO_M1_d N_net_m1_VDDO_res_M1_g N_U14_pgate_tol_M1_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M41 N_U14_padr_M41_d N_net_m41_VSSO_res_M41_g N_VSSO_M41_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U14_padr_M41@2_d N_net_m41_VSSO_res_M41@2_g N_VSSO_M41_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U9_U33_source_M39_d N_U14_padr_M39_g N_VSSO_M39_s N_VSS_M3_b NHV
+ L=3.6e-07 W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M40 N_U9_U41_gate_M40_d N_U14_padr_M40_g N_U9_U33_source_M39_d N_VSS_M3_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M38 N_VDDO_M38_d N_U9_U41_gate_M38_g N_U9_U33_source_M38_s N_VSS_M3_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M42 N_U9_U43_drain_M42_d N_U9_U41_gate_M42_g N_VSSO_M42_s N_VSS_M3_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M42@2 N_U9_U43_drain_M42_d N_U9_U41_gate_M42@2_g N_VSSO_M42@2_s N_VSS_M3_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M43 N_CIN_M43_d N_U9_U43_drain_M43_g N_VSS_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M4 N_U14_pgate_tol_M4_s N_net_m4_VSSO_res_M4_g N_U14_pgate_tol_M4_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VSSO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VSSO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VDDO_M4_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_U14_pgate_tol_M2_d N_net_m2_VSSO_res_M2_g N_VDDO_M2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M35 N_U14_padr_M35_d N_net_m35_VDDO_res_M35_g N_VDDO_M35_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U14_padr_M35_d N_net_m35_VDDO_res_M35@2_g N_VDDO_M35@2_s N_VDDO_M4_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M34 N_U9_U41_source_M34_d N_U14_padr_M34_g N_VDDO_M34_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M33 N_U9_U41_gate_M33_d N_U14_padr_M33_g N_U9_U41_source_M34_d N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M32 N_VSSO_M32_d N_U9_U41_gate_M32_g N_U9_U41_source_M32_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M36 N_U9_U43_drain_M36_d N_U9_U41_gate_M36_g N_VDDO_M36_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M36@2 N_U9_U43_drain_M36_d N_U9_U41_gate_M36@2_g N_VDDO_M36@2_s N_VDDO_M4_b PHV
+ L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M37 N_CIN_M37_d N_U9_U43_drain_M37_g N_VDD_M37_s N_VDD_M37_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M37@2 N_CIN_M37@2_d N_U9_U43_drain_M37@2_g N_VDD_M37_s N_VDD_M37_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M37@3 N_CIN_M37@2_d N_U9_U43_drain_M37@3_g N_VDD_M37@3_s N_VDD_M37_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M37@4 N_CIN_M37@4_d N_U9_U43_drain_M37@4_g N_VDD_M37@3_s N_VDD_M37_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM35 N_net_m35_VDDO_res_RM35_pos N_VDDO_RM35_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_VDDO_RM3_pos N_net_m3_VDDO_res_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM1 N_VDDO_RM1_pos N_net_m1_VDDO_res_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_net_m2_VSSO_res_RM2_pos N_VSSO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM41 N_VSSO_RM41_pos N_net_m41_VSSO_res_RM41_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d31.dist.sp.PC3D31.pxi"
*
.ends
*
*
* File: pc3d31u.dist.sp
* Created: Sun Jul  4 12:35:36 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3d31u.dist.sp.pex"
.subckt pc3d31u  CIN PAD VDD VSS VDDO VSSO 
* 
M8 N_PAD_M14_d N_U14_MN4$11_gate_M8_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M15_d N_U14_MN4$11_gate_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M16_d N_U14_MN4$11_gate_M10_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U14_MN4$11_gate_M11_g N_VSSO_M8_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M18_d N_U14_MN4$11_gate_M12_g N_VSSO_M12_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M19_d N_U14_MN4$11_gate_M13_g N_VSSO_M10_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U14_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M5_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR20 N_U14_MN4$11_gate_R20_pos N_VSSO_R20_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M14 N_PAD_M14_d N_U14_MN4$11_gate_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_U14_MN4$11_gate_M15_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U14_MN4$11_gate_M16_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U14_MN4$11_gate_M17_g N_VSSO_M16_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U14_MN4$11_gate_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M19_d N_U14_MN4$11_gate_M19_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
M21 N_VDDO_M21_d N_U14_pgate_tol_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M22 N_VDDO_M25_d N_U14_pgate_tol_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_U14_pgate_tol_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U14_pgate_tol_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U14_pgate_tol_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U14_pgate_tol_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U14_pgate_tol_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U14_pgate_tol_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U14_pgate_tol_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U14_pgate_tol_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U14_pgate_tol_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U14_pgate_tol_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR6 N_X26/noxref_9_R6_pos N_PAD_R6_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR7 N_X26/noxref_9_R7_pos N_U14_padr_R7_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M4 N_U14_pgate_tol_M4_s N_net_m4_VDDO_res_M4_g N_U14_pgate_tol_M4_s N_VSS_M4_b
+ NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M4@2 N_U14_pgate_tol_M4@2_s N_net_m4_VDDO_res_M4@2_g N_U14_pgate_tol_M4@2_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M4@3 N_U14_pgate_tol_M4@3_s N_net_m4_VDDO_res_M4@3_g N_U14_pgate_tol_M4@3_s
+ N_VSS_M4_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M2 N_VDDO_M2_d N_net_m2_VDDO_res_M2_g N_U14_pgate_tol_M2_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U14_padr_M42_d N_net_m42_VSSO_res_M42_g N_VSSO_M42_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M42@2 N_U14_padr_M42@2_d N_net_m42_VSSO_res_M42@2_g N_VSSO_M42_s N_VSS_M4_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40 N_U9_U33_source_M40_d N_U14_padr_M40_g N_VSSO_M40_s N_VSS_M4_b NHV
+ L=3.6e-07 W=9.5e-06 AD=4.34548e-12 AS=5.89e-12 PD=1.26503e-05 PS=2.024e-05
M41 N_U9_U41_gate_M41_d N_U14_padr_M41_g N_U9_U33_source_M40_d N_VSS_M4_b NHV
+ L=3.6e-07 W=6e-06 AD=3.9e-12 AS=2.74452e-12 PD=1.33e-05 PS=7.98968e-06
M39 N_VDDO_M39_d N_U9_U41_gate_M39_g N_U9_U33_source_M39_s N_VSS_M4_b NHV
+ L=3.6e-07 W=2.5e-06 AD=1.55e-12 AS=1.55e-12 PD=6.24e-06 PS=6.24e-06
M43 N_U9_U43_drain_M43_d N_U9_U41_gate_M43_g N_VSSO_M43_s N_VSS_M4_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M43@2 N_U9_U43_drain_M43_d N_U9_U41_gate_M43@2_g N_VSSO_M43@2_s N_VSS_M4_b NHV
+ L=3.6e-07 W=7.5e-06 AD=3.075e-12 AS=4.65e-12 PD=8.32e-06 PS=1.624e-05
M44 N_CIN_M44_d N_U9_U43_drain_M44_g N_VSS_M44_s N_VSS_M4_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M5 N_U14_pgate_tol_M5_s N_net_m5_VSSO_res_M5_g N_U14_pgate_tol_M5_s N_VDDO_M5_b
+ PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M5@2 N_U14_pgate_tol_M5@2_s N_net_m5_VSSO_res_M5@2_g N_U14_pgate_tol_M5@2_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M5@3 N_U14_pgate_tol_M5@3_s N_net_m5_VSSO_res_M5@3_g N_U14_pgate_tol_M5@3_s
+ N_VDDO_M5_b PHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M3 N_U14_pgate_tol_M3_d N_net_m3_VSSO_res_M3_g N_VDDO_M3_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M36 N_U14_padr_M36_d N_net_m36_VDDO_res_M36_g N_VDDO_M36_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M36@2 N_U14_padr_M36_d N_net_m36_VDDO_res_M36@2_g N_VDDO_M36@2_s N_VDDO_M5_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35 N_U9_U41_source_M35_d N_U14_padr_M35_g N_VDDO_M35_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=1.1e-05 AD=4.51e-12 AS=6.82e-12 PD=1.182e-05 PS=2.324e-05
M34 N_U9_U41_gate_M34_d N_U14_padr_M34_g N_U9_U41_source_M35_d N_VDDO_M5_b PHV
+ L=3.6e-07 W=1.1e-05 AD=6.82e-12 AS=4.51e-12 PD=2.324e-05 PS=1.182e-05
M33 N_VSSO_M33_d N_U9_U41_gate_M33_g N_U9_U41_source_M33_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=4.96e-12 PD=1.724e-05 PS=1.724e-05
M37 N_U9_U43_drain_M37_d N_U9_U41_gate_M37_g N_VDDO_M37_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=2e-05 AD=8.48e-12 AS=1.24e-11 PD=2.2208e-05 PS=4.124e-05
M37@2 N_U9_U43_drain_M37_d N_U9_U41_gate_M37@2_g N_VDDO_M37@2_s N_VDDO_M5_b PHV
+ L=3.6e-07 W=1.75e-05 AD=7.42e-12 AS=1.085e-11 PD=1.9432e-05 PS=3.624e-05
M38 N_CIN_M38_d N_U9_U43_drain_M38_g N_VDD_M38_s N_VDD_M38_b PHV L=3.6e-07
+ W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
M38@2 N_CIN_M38@2_d N_U9_U43_drain_M38@2_g N_VDD_M38_s N_VDD_M38_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M38@3 N_CIN_M38@2_d N_U9_U43_drain_M38@3_g N_VDD_M38@3_s N_VDD_M38_b PHV
+ L=3.6e-07 W=9e-06 AD=3.69e-12 AS=3.69e-12 PD=9.82e-06 PS=9.82e-06
M38@4 N_CIN_M38@4_d N_U9_U43_drain_M38@4_g N_VDD_M38@3_s N_VDD_M38_b PHV
+ L=3.6e-07 W=9e-06 AD=5.58e-12 AS=3.69e-12 PD=1.924e-05 PS=9.82e-06
XRM36 N_net_m36_VDDO_res_RM36_pos N_VDDO_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM5 N_VSSO_RM5_pos N_net_m5_VSSO_res_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM4 N_VDDO_RM4_pos N_net_m4_VDDO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM2 N_VDDO_RM2_pos N_net_m2_VDDO_res_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM3 N_net_m3_VSSO_res_RM3_pos N_VSSO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM42 N_VSSO_RM42_pos N_net_m42_VSSO_res_RM42_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
*
.include "pc3d31u.dist.sp.PC3D31U.pxi"
*
.ends
*
*
* File: pc3o01hv.dist.sp
* Created: Sun Jul  4 12:37:32 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o01hv.dist.sp.pex"
.subckt pc3o01hv  PAD I VDD VSS VDDO VSSO 
* 
M17 N_PAD_M23_d N_U29_U74$9_gate_M17_g N_VSSO_M17_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M24_d N_U29_U74$9_gate_M18_g N_VSSO_M18_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M19 N_PAD_M25_d N_U29_U74$9_gate_M19_g N_VSSO_M19_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M26_d N_U29_U74$9_gate_M20_g N_VSSO_M17_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M21 N_PAD_M15_d N_U29_U74$9_gate_M21_g N_VSSO_M21_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M22 N_PAD_M16_d N_U29_U74$9_gate_M22_g N_VSSO_M19_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR39 N_VSSO_R39_pos N_U29_U74$9_gate_R39_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR40 N_U29_U37_r2_R40_pos N_VDDO_R40_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M23 N_PAD_M23_d N_U29_U74$9_gate_M23_g N_VSSO_M23_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M24_d N_U29_U74$9_gate_M24_g N_VSSO_M23_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M25_d N_U29_U74$9_gate_M25_g N_VSSO_M25_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M26_d N_U29_U74$9_gate_M26_g N_VSSO_M25_s N_VSSO_M23_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M15_d N_ngate_M15_g N_VSSO_M15_s N_VSSO_M23_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_ngate_M16_g N_VSSO_M15_s N_VSSO_M23_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR13 U29_U69_padr N_noxref_2_R13_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR14 N_noxref_2_R14_pos N_PAD_R14_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M29 N_VDDO_M29_d N_U29_U37_r2_M29_g N_PAD_M29_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M30 N_VDDO_M31_d N_U29_U37_r2_M30_g N_PAD_M29_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M38_d N_pgate_M27_g N_PAD_M27_s N_VDDO_M31_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_pgate_M28_g N_PAD_M27_s N_VDDO_M31_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M31 N_VDDO_M31_d N_U29_U37_r2_M31_g N_PAD_M31_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U37_r2_M32_g N_PAD_M31_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U37_r2_M33_g N_PAD_M33_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U37_r2_M34_g N_PAD_M33_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_VDDO_M34_d N_U29_U37_r2_M35_g N_PAD_M35_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U29_U37_r2_M36_g N_PAD_M35_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M37 N_VDDO_M36_d N_U29_U37_r2_M37_g N_PAD_M37_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M38 N_VDDO_M38_d N_U29_U37_r2_M38_g N_PAD_M37_s N_VDDO_M31_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M1 N_ngate_M1_d N_U28_ISHF_M1_g N_VSSO_M1_s N_VSS_M1_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M1@2 N_ngate_M1_d N_U28_ISHF_M1@2_g N_VSSO_M1@2_s N_VSS_M1_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M2 N_pgate_M2_d N_net_m2_VDDO_res_M2_g N_ngate_M2_s N_VSS_M1_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M2@2 N_pgate_M2@2_d N_net_m2_VDDO_res_M2@2_g N_ngate_M2_s N_VSS_M1_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M2@3 N_pgate_M2@2_d N_net_m2_VDDO_res_M2@3_g N_ngate_M2@3_s N_VSS_M1_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9 N_U28_U13_MPLL1_dr_M9_d N_I_M9_g N_VSSO_M9_s N_VSS_M1_b NHV L=3.6e-07
+ W=8e-06 AD=4.96e-12 AS=5.12e-12 PD=1.724e-05 PS=1.728e-05
M10 N_U28_ISHF_M10_d N_U28_U13_MPLL1_dr_M10_g N_VSSO_M10_s N_VSS_M1_b NHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M10@2 N_U28_ISHF_M10_d N_U28_U13_MPLL1_dr_M10@2_g N_VSSO_M10@2_s N_VSS_M1_b NHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@3 N_U28_ISHF_M10@3_d N_U28_U13_MPLL1_dr_M10@3_g N_VSSO_M10@2_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@4 N_U28_ISHF_M10@3_d N_U28_U13_MPLL1_dr_M10@4_g N_VSSO_M10@4_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@5 N_U28_ISHF_M10@5_d N_U28_U13_MPLL1_dr_M10@5_g N_VSSO_M10@4_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M10@6 N_U28_ISHF_M10@5_d N_U28_U13_MPLL1_dr_M10@6_g N_VSSO_M10@6_s N_VSS_M1_b
+ NHV L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M5 N_U28_U13_U6_drain_M5_d N_net_m5_VSS_res_M5_g N_VSS_M5_s N_VSS_M1_b N18
+ L=1.8e-07 W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M3 N_pgate_M3_d N_U28_ISHF_M3_g N_VDDO_M3_s N_VDDO_M3_b PHV L=3.6e-07 W=2e-05
+ AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M3@2 N_pgate_M3@2_d N_U28_ISHF_M3@2_g N_VDDO_M3_s N_VDDO_M3_b PHV L=3.6e-07
+ W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M4 N_ngate_M4_d N_net_m4_VSSO_res_M4_g N_pgate_M4_s N_VDDO_M3_b PHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M4@2 N_ngate_M4_d N_net_m4_VSSO_res_M4@2_g N_pgate_M4@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M4@3 N_ngate_M4@3_d N_net_m4_VSSO_res_M4@3_g N_pgate_M4@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7 N_U28_U13_MPLL1_dr_M7_d N_I_M7_g N_VDDO_M7_s N_VDDO_M3_b PHV L=3.6e-07
+ W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M8 N_U28_ISHF_M8_d N_U28_U13_MPLL1_dr_M8_g N_VDDO_M8_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M8@2 N_U28_ISHF_M8_d N_U28_U13_MPLL1_dr_M8@2_g N_VDDO_M8@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@3 N_U28_ISHF_M8@3_d N_U28_U13_MPLL1_dr_M8@3_g N_VDDO_M8@2_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@4 N_U28_ISHF_M8@3_d N_U28_U13_MPLL1_dr_M8@4_g N_VDDO_M8@4_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@5 N_U28_ISHF_M8@5_d N_U28_U13_MPLL1_dr_M8@5_g N_VDDO_M8@4_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=2.46e-12 PD=6.82e-06 PS=6.82e-06
M8@6 N_U28_ISHF_M8@5_d N_U28_U13_MPLL1_dr_M8@6_g N_VDDO_M8@6_s N_VDDO_M3_b PHV
+ L=3.6e-07 W=6e-06 AD=2.46e-12 AS=3.72e-12 PD=6.82e-06 PS=1.324e-05
M6 N_U28_U13_U6_drain_M6_d N_net_m6_VDD_res_M6_g N_VDD_M6_s N_VDD_M6_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M6@2 N_U28_U13_U6_drain_M6_d N_net_m6_VDD_res_M6@2_g N_VDD_M6@2_s N_VDD_M6_b
+ P18 L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D12 N_VSS_M1_b N_I_D12_neg DN18  AREA=1e-12 PJ=4e-06
XRM2 N_net_m2_VDDO_res_RM2_pos N_VDDO_RM2_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM4 N_net_m4_VSSO_res_RM4_pos N_VSSO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM5 N_net_m5_VSS_res_RM5_pos N_VSS_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM6 N_net_m6_VDD_res_RM6_pos N_VDD_RM6_neg RPMPOLY2T w=2e-06 l=6.455e-06 
c_1 U29_U69_padr 0 17.4974f
*
.include "pc3o01hv.dist.sp.PC3O01HV.pxi"
*
.ends
*
*
* File: pc3o01.dist.sp
* Created: Sun Jul  4 12:35:39 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o01.dist.sp.pex"
.subckt pc3o01  PAD I VDD VSS VDDO VSSO 
* 
M29 N_ngate_M29_d N_U28_ISHF_M29_g N_VSSO_M29_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M29@2 N_ngate_M29_d N_U28_ISHF_M29@2_g N_VSSO_M29@2_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M30 N_pgate_M30_d N_net_m30_VDDO_res_M30_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M30@2 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@2_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M30@3 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@3_g N_ngate_M30@3_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_VDDO_M37_d N_U28_U16_MN1_drai_M37_g N_U28_U16_MPLL1_dr_M37_s N_VSS_M29_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M35 N_U28_U16_MPLL1_dr_M35_d N_I_M35_g N_VSSO_M35_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M35@2 N_U28_U16_MPLL1_dr_M35@2_d N_I_M35@2_g N_VSSO_M35_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36 N_U28_ISHF_M36_d N_U28_U16_MN1_drai_M36_g N_VSSO_M36_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36@2 N_U28_ISHF_M36@2_d N_U28_U16_MN1_drai_M36@2_g N_VSSO_M36_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_PAD_M11_d N_U29_U74$9_gate_M5_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M12_d N_U29_U74$9_gate_M6_g N_VSSO_M6_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M13_d N_U29_U74$9_gate_M7_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U29_U74$9_gate_M8_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M3_d N_U29_U74$9_gate_M9_g N_VSSO_M9_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M4_d N_U29_U74$9_gate_M10_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_U28_U16_MN1_drai_M38_d N_I_M38_g N_VSS_M38_s N_VSS_M29_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M31 N_pgate_M31_d N_U28_ISHF_M31_g N_VDDO_M31_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M31@2 N_pgate_M31@2_d N_U28_ISHF_M31@2_g N_VDDO_M31_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M32 N_ngate_M32_d N_net_m32_VSSO_res_M32_g N_pgate_M32_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_ngate_M32_d N_net_m32_VSSO_res_M32@2_g N_pgate_M32@2_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M32@3 N_ngate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_pgate_M32@2_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33 N_U28_U16_MPLL1_dr_M33_d N_U28_ISHF_M33_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M34 N_U28_ISHF_M34_d N_U28_U16_MPLL1_dr_M34_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M39 N_U28_U16_MN1_drai_M39_d N_I_M39_g N_VDD_M39_s N_VDD_M39_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M39@2 N_U28_U16_MN1_drai_M39_d N_I_M39@2_g N_VDD_M39@2_s N_VDD_M39_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D40 N_VSS_M29_b N_I_D40_neg DN18  AREA=2.5e-13 PJ=2e-06
XR27 N_VSSO_R27_pos N_U29_U74$9_gate_R27_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR28 N_U29_U37_r2_R28_pos N_VDDO_R28_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M11 N_PAD_M11_d N_U29_U74$9_gate_M11_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_U74$9_gate_M12_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U74$9_gate_M13_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U29_U74$9_gate_M14_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M3 N_PAD_M3_d N_ngate_M3_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_ngate_M4_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR1 U29_U69_padr N_noxref_11_R1_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR2 N_noxref_11_R2_pos N_PAD_R2_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XRM30 N_net_m30_VDDO_res_RM30_pos N_VDDO_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M17 N_VDDO_M17_d N_U29_U37_r2_M17_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M18 N_VDDO_M19_d N_U29_U37_r2_M18_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M15 N_VDDO_M26_d N_pgate_M15_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M16 N_VDDO_M16_d N_pgate_M16_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M19 N_VDDO_M19_d N_U29_U37_r2_M19_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U29_U37_r2_M20_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U29_U37_r2_M21_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U29_U37_r2_M22_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U29_U37_r2_M23_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U29_U37_r2_M24_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M24_d N_U29_U37_r2_M25_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U37_r2_M26_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U29_U69_padr 0 17.4974f
*
.include "pc3o01.dist.sp.PC3O01.pxi"
*
.ends
*
*
* File: pc3o02.dist.sp
* Created: Sun Jul  4 12:37:43 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o02.dist.sp.pex"
.subckt pc3o02  PAD I VDD VSS VDDO VSSO 
* 
M23 N_PAD_M27_d N_U29_U74$7_gate_M23_g N_VSSO_M23_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M24 N_PAD_M28_d N_U29_U74$7_gate_M24_g N_VSSO_M24_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M21 N_PAD_M29_d N_ngate_M21_g N_VSSO_M21_s N_VSSO_M27_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M25 N_PAD_M30_d N_U29_U74$7_gate_M25_g N_VSSO_M23_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_PAD_M19_d N_U29_U74$7_gate_M26_g N_VSSO_M26_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M22 N_PAD_M20_d N_ngate_M22_g N_VSSO_M21_s N_VSSO_M27_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR45 N_VSSO_R45_pos N_U29_U74$7_gate_R45_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR46 N_U29_U37_r2_R46_pos N_VDDO_R46_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M27 N_PAD_M27_d N_U29_U74$7_gate_M27_g N_VSSO_M27_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M28 N_PAD_M28_d N_U29_U74$7_gate_M28_g N_VSSO_M27_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M29 N_PAD_M29_d N_U29_U74$7_gate_M29_g N_VSSO_M29_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M30 N_PAD_M30_d N_U29_U74$7_gate_M30_g N_VSSO_M29_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M19 N_PAD_M19_d N_U30_ngate2_M19_g N_VSSO_M19_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_PAD_M20_d N_U30_ngate2_M20_g N_VSSO_M19_s N_VSSO_M27_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR31 U29_U69_padr N_noxref_2_R31_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR32 N_noxref_2_R32_pos N_PAD_R32_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M37 N_VDDO_M37_d N_U29_U37_r2_M37_g N_PAD_M37_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M38 N_VDDO_M39_d N_U29_U37_r2_M38_g N_PAD_M37_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M36_d N_pgate_M33_g N_PAD_M33_s N_VDDO_M39_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_pgate_M34_g N_PAD_M33_s N_VDDO_M39_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M39 N_VDDO_M39_d N_U29_U37_r2_M39_g N_PAD_M39_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M40 N_VDDO_M40_d N_U29_U37_r2_M40_g N_PAD_M39_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M41 N_VDDO_M40_d N_U29_U37_r2_M41_g N_PAD_M41_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M42 N_VDDO_M42_d N_U29_U37_r2_M42_g N_PAD_M41_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M42_d N_U29_U37_r2_M43_g N_PAD_M43_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M44 N_VDDO_M44_d N_U29_U37_r2_M44_g N_PAD_M43_s N_VDDO_M39_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M35 N_VDDO_M44_d N_pgate_M35_g N_PAD_M35_s N_VDDO_M39_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_pgate_M36_g N_PAD_M35_s N_VDDO_M39_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_ngate_M7_d N_U28_ISHF_M7_g N_VSSO_M7_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M7@2 N_ngate_M7_d N_U28_ISHF_M7@2_g N_VSSO_M7@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M8 N_pgate_M8_d N_net_m8_VDDO_res_M8_g N_ngate_M8_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_pgate_M8@2_d N_net_m8_VDDO_res_M8@2_g N_ngate_M8_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_pgate_M8@2_d N_net_m8_VDDO_res_M8@3_g N_ngate_M8@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M15 N_VDDO_M15_d N_U28_U16_MN1_drai_M15_g N_U28_U16_MPLL1_dr_M15_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U28_U16_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U28_U16_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U28_ISHF_M14_d N_U28_U16_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U28_ISHF_M14@2_d N_U28_U16_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U28_U16_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M9 N_pgate_M9_d N_U28_ISHF_M9_g N_VDDO_M9_s N_VDDO_M6_b PHV L=3.6e-07 W=2e-05
+ AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M9@2 N_pgate_M9@2_d N_U28_ISHF_M9@2_g N_VDDO_M9_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M10 N_ngate_M10_d N_net_m10_VSSO_res_M10_g N_pgate_M10_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M10@2 N_ngate_M10_d N_net_m10_VSSO_res_M10@2_g N_pgate_M10@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M10@3 N_ngate_M10@3_d N_net_m10_VSSO_res_M10@3_g N_pgate_M10@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M11 N_U28_U16_MPLL1_dr_M11_d N_U28_ISHF_M11_g N_VDDO_M11_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U28_ISHF_M12_d N_U28_U16_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M17 N_U28_U16_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U28_U16_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D18 N_VSS_M3_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM8 N_net_m8_VDDO_res_RM8_pos N_VDDO_RM8_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM10 N_net_m10_VSSO_res_RM10_pos N_VSSO_RM10_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.5032f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pc3o02.dist.sp.PC3O02.pxi"
*
.ends
*
*
* File: pc3o03.dist.sp
* Created: Sun Jul  4 12:38:48 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o03.dist.sp.pex"
.subckt pc3o03  PAD I VDD VSS VDDO VSSO 
* 
M13 N_PAD_M17_d N_U29_U76_r1_M13_g N_VSSO_M13_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M18_d N_U29_U76_r1_M14_g N_VSSO_M14_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M7_d N_U30_ngate2_M9_g N_VSSO_M9_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M8_d N_U29_U76_r1_M15_g N_VSSO_M13_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M11_d N_U29_U76_r1_M16_g N_VSSO_M16_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M12_d N_U30_ngate2_M10_g N_VSSO_M9_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M17 N_PAD_M17_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U29_U76_r1_M18_g N_VSSO_M17_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M7_d N_ngate_M7_g N_VSSO_M7_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_ngate_M8_g N_VSSO_M7_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U29_ngate3_M11_g N_VSSO_M11_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_ngate3_M12_g N_VSSO_M11_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR31 U29_U69_padr N_noxref_2_R31_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR32 N_noxref_2_R32_pos N_PAD_R32_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U29_U37_r2_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U29_U37_r2_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U37_r2_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U37_r2_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U37_r2_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U37_r2_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U29_ngate3_M34_d N_U30_ngatex_M34_g N_VSSO_M34_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U28_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U28_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U28_U13_MN1_drai_M45_g N_U28_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U28_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U28_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U28_ISHF_M44_d N_U28_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U28_ISHF_M44@2_d N_U28_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U28_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M33 N_U29_ngate3_M33_d N_U30_ngatex_M33_g N_U30_ngate2_M33_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U28_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U28_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U28_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U28_U13_MPLL1_dr_M41_d N_U28_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U28_ISHF_M42_d N_U28_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U28_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U28_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.5122f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pc3o03.dist.sp.PC3O03.pxi"
*
.ends
*
*
* File: pc3o04.dist.sp
* Created: Sun Jul  4 12:38:52 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o04.dist.sp.pex"
.subckt pc3o04  PAD I VDD VSS VDDO VSSO 
* 
M15 N_PAD_M8_d N_U29_U76_r1_M15_g N_VSSO_M15_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M9_d N_ngate_M7_g N_VSSO_M7_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M17_d N_U29_ngate3_M13_g N_VSSO_M13_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U29_U76_r1_M16_g N_VSSO_M15_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U30_ngate2_M10_g N_VSSO_M10_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M14 N_PAD_M12_d N_U29_ngate3_M14_g N_VSSO_M13_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M8 N_PAD_M8_d N_ngate_M8_g N_VSSO_M8_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M9_d N_ngate_M9_g N_VSSO_M8_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U29_U76_r1_M18_g N_VSSO_M17_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U30_ngate2_M11_g N_VSSO_M11_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U30_ngate2_M12_g N_VSSO_M11_s N_VSSO_M8_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR31 U29_U69_padr N_noxref_2_R31_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR32 N_noxref_2_R32_pos N_PAD_R32_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M27 N_VDDO_M27_d N_U29_U37_r2_M27_g N_PAD_M27_s N_VDDO_M29_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M28 N_VDDO_M29_d N_U29_U37_r2_M28_g N_PAD_M27_s N_VDDO_M29_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M26_d N_pgate_M19_g N_PAD_M19_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_pgate_M20_g N_PAD_M19_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M29 N_VDDO_M29_d N_U29_U37_r2_M29_g N_PAD_M29_s N_VDDO_M29_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U37_r2_M30_g N_PAD_M29_s N_VDDO_M29_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_pgate_M21_g N_PAD_M21_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_pgate_M22_g N_PAD_M21_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M24_d N_pgate_M25_g N_PAD_M25_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_pgate_M26_g N_PAD_M25_s N_VDDO_M29_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U29_ngate3_M34_d N_U30_ngatex_M34_g N_VSSO_M34_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U28_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U28_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U28_U13_MN1_drai_M45_g N_U28_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U28_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U28_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U28_ISHF_M44_d N_U28_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U28_ISHF_M44@2_d N_U28_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U28_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M33 N_U29_ngate3_M33_d N_U30_ngatex_M33_g N_U30_ngate2_M33_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U28_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U28_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U28_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U28_U13_MPLL1_dr_M41_d N_U28_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U28_ISHF_M42_d N_U28_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U28_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U28_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.4923f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pc3o04.dist.sp.PC3O04.pxi"
*
.ends
*
*
* File: pc3o05.dist.sp
* Created: Sun Jul  4 12:40:47 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3o05.dist.sp.pex"
.subckt pc3o05  PAD I VDD VSS VDDO VSSO 
* 
M13 N_PAD_M15_d N_ngate_M13_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M16_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M9_d N_U30_ngate2_M7_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M10_d N_ngate_M14_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M11_d N_U29_U76_r1_M18_g N_VSSO_M18_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M12_d N_U30_ngate2_M8_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M15 N_PAD_M15_d N_ngate_M15_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_ngate_M16_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M9_d N_U30_ngate2_M9_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U30_ngate2_M10_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U29_ngate3_M11_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_ngate3_M12_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 U29_U69_padr N_noxref_2_R19_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR20 N_noxref_2_R20_pos N_PAD_R20_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M33 N_VDDO_M33_d N_U29_U37_r2_M33_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M25_d N_U29_U37_r2_M34_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_pgate_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_pgate_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_pgate_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_pgate_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_pgate_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_pgate_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_pgate_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_pgate_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M22 N_U29_ngate3_M22_d N_U30_ngatex_M22_g N_VSSO_M22_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U27_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U27_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U27_U13_MN1_drai_M45_g N_U27_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U27_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U27_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U27_ISHF_M44_d N_U27_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U27_ISHF_M44@2_d N_U27_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U27_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M21 N_U29_ngate3_M21_d N_U30_ngatex_M21_g N_U30_ngate2_M21_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U27_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U27_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U27_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U27_U13_MPLL1_dr_M41_d N_U27_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U27_ISHF_M42_d N_U27_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U27_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U27_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.4884f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pc3o05.dist.sp.PC3O05.pxi"
*
.ends
*
*
* File: pc3t01d.dist.sp
* Created: Sun Jul  4 12:42:11 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t01d.dist.sp.pex"
.subckt pc3t01d  PAD I OEN VDD VSS VDDO VSSO 
* 
M56 N_U27_padr_M56_d N_net_m56_VDDO_res_M56_g U28_U22_source N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M57 U28_U22_source N_net_m57_VDDO_res_M57_g N_VSSO_M57_s N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM56 N_net_m56_VDDO_res_RM56_pos N_VDDO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM57 N_VDDO_RM56_neg N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M61 N_U27_padr_M61_d N_net_m61_VSSO_res_M61_g N_VSSO_M61_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M61@2 N_U27_padr_M61@2_d N_net_m61_VSSO_res_M61@2_g N_VSSO_M61_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62 N_U29_MPI1_drain_M62_d N_U27_padr_M62_g N_VSSO_M62_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M60 N_U27_padr_M60_d N_net_m60_VDDO_res_M60_g N_VDDO_M60_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 U29_MPI2_drain N_U27_padr_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M59 N_U29_MPI1_drain_M59_d N_U27_padr_M59_g U29_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM60 N_net_m60_VDDO_res_RM60_pos N_VDDO_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM61 N_VSSO_RM61_pos N_net_m61_VSSO_res_RM61_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_MPI2_drain 0 0.0289375f
*
.include "pc3t01d.dist.sp.PC3T01D.pxi"
*
.ends
*
*
* File: pc3t01.dist.sp
* Created: Sun Jul  4 12:40:31 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t01.dist.sp.pex"
.subckt pc3t01  PAD I OEN VDD VSS VDDO VSSO 
* 
M32 N_PAD_M33_d N_U27_U69$9_gate_M32_g N_VSSO_M32_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M33_d N_U27_U69$9_gate_M33_g N_VSSO_M33_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M35_d N_U27_U69$9_gate_M34_g N_VSSO_M34_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M35_d N_U27_U69$9_gate_M35_g N_VSSO_M32_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M37_d N_U27_U69$9_gate_M36_g N_VSSO_M36_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M37 N_PAD_M37_d N_U27_U69$9_gate_M37_g N_VSSO_M34_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M39_d N_U27_U69$9_gate_M38_g N_VSSO_M38_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M39 N_PAD_M39_d N_U27_U69$9_gate_M39_g N_VSSO_M36_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M30 N_PAD_M40_d N_U15_ngate_M30_g N_VSSO_M30_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U27_U69$9_gate_M40_g N_VSSO_M38_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M31_d N_U27_U69$9_gate_M41_g N_VSSO_M41_s N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M31 N_PAD_M31_d N_U15_ngate_M31_g N_VSSO_M30_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M55 N_U15_pgate_M55_d N_net_m55_VSSO_res_M55_g N_U27_U72_pgate_M55_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M55@2 N_U15_pgate_M55_d N_net_m55_VSSO_res_M55@2_g N_U27_U72_pgate_M55@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@3 N_U15_pgate_M55@3_d N_net_m55_VSSO_res_M55@3_g N_U27_U72_pgate_M55@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@4 N_U15_pgate_M55@3_d N_net_m55_VSSO_res_M55@4_g N_U27_U72_pgate_M55@4_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M55@5 N_U15_pgate_M55@5_d N_net_m55_VSSO_res_M55@5_g N_U27_U72_pgate_M55@4_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR58 N_U27_U69$9_gate_R58_pos N_VSSO_R58_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR56 N_noxref_2_R56_pos N_PAD_R56_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR57 N_noxref_2_R57_pos N_U27_padr_R57_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M44 N_VDDO_M44_d N_U27_U71_UN_P_TOP_M44_g N_PAD_M44_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M45 N_VDDO_M46_d N_U27_U71_UN_P_TOP_M45_g N_PAD_M44_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M42 N_VDDO_M53_d N_U27_U72_pgate_M42_g N_PAD_M42_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M43_d N_U27_U72_pgate_M43_g N_PAD_M42_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M46 N_VDDO_M46_d N_U27_U71_UN_P_TOP_M46_g N_PAD_M46_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M47 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M47_g N_PAD_M46_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M48 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M48_g N_PAD_M48_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M49 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M49_g N_PAD_M48_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M50_g N_PAD_M50_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M51 N_VDDO_M51_d N_U27_U71_UN_P_TOP_M51_g N_PAD_M50_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M51_d N_U27_U71_UN_P_TOP_M52_g N_PAD_M52_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M53_d N_U27_U71_UN_P_TOP_M53_g N_PAD_M52_s N_VDDO_M46_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_U15_pgate_M54_d N_net_m54_VDDO_res_M54_g N_U27_U72_pgate_M54_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M54@2 N_U15_pgate_M54_d N_net_m54_VDDO_res_M54@2_g N_U27_U72_pgate_M54@2_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M54@3 N_U15_pgate_M54@3_d N_net_m54_VDDO_res_M54@3_g N_U27_U72_pgate_M54@2_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M59 N_VDDO_M59_d N_net_m59_VDDO_res_M59_g N_U27_U71_UN_P_TOP_M59_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M4 N_U27_padr_M4_d N_net_m4_VSSO_res_M4_g N_VSSO_M4_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M4@2 N_U27_padr_M4@2_d N_net_m4_VSSO_res_M4@2_g N_VSSO_M4_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_U28_MPI1_drain_M5_d N_U27_padr_M5_g N_VSSO_M5_s N_VSS_M54_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M27 N_U15_U12_oenb_M27_d N_U15_U15_OUTSHIFT_M27_g N_VSSO_M27_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M6 N_U15_ngate_M6_d N_U15_ISHF_M6_g N_VSSO_M6_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M6@2 N_U15_ngate_M6_d N_U15_ISHF_M6@2_g N_VSSO_M6@2_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M26 N_U15_ngate_M26_d N_U15_U15_OUTSHIFT_M26_g N_VSSO_M6@2_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M7 N_U15_pgate_M7_d N_U15_U12_oenb_M7_g N_U15_ngate_M7_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7@2 N_U15_pgate_M7@2_d N_U15_U12_oenb_M7@2_g N_U15_ngate_M7_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M7@3 N_U15_pgate_M7@2_d N_U15_U12_oenb_M7@3_g N_U15_ngate_M7@3_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M20 N_U15_U15_MPLL1_dr_M20_d N_OEN_M20_g N_VSSO_M20_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M22 N_VDDO_M22_d N_U15_U15_MN1_drai_M22_g N_U15_U15_MPLL1_dr_M22_s N_VSS_M54_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M20@2 N_U15_U15_MPLL1_dr_M20@2_d N_OEN_M20@2_g N_VSSO_M20_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M21 N_U15_U15_OUTSHIFT_M21_d N_U15_U15_MN1_drai_M21_g N_VSSO_M21_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M21@2 N_U15_U15_OUTSHIFT_M21@2_d N_U15_U15_MN1_drai_M21@2_g N_VSSO_M21_s
+ N_VSS_M54_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M14 N_VDDO_M14_d N_U15_U14_MN1_drai_M14_g N_U15_U14_MPLL1_dr_M14_s N_VSS_M54_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M12 N_U15_U14_MPLL1_dr_M12_d N_I_M12_g N_VSSO_M12_s N_VSS_M54_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M12@2 N_U15_U14_MPLL1_dr_M12@2_d N_I_M12@2_g N_VSSO_M12_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13 N_U15_ISHF_M13_d N_U15_U14_MN1_drai_M13_g N_VSSO_M13_s N_VSS_M54_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U15_ISHF_M13@2_d N_U15_U14_MN1_drai_M13@2_g N_VSSO_M13_s N_VSS_M54_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M15 N_U15_U14_MN1_drai_M15_d N_I_M15_g N_VSS_M15_s N_VSS_M54_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M23 N_U15_U15_MN1_drai_M23_d N_OEN_M23_g N_VSS_M15_s N_VSS_M54_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M60 N_U27_U71_UN_P_TOP_M60_d N_net_m60_VSSO_res_M60_g N_VDDO_M60_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M3 N_U27_padr_M3_d N_net_m3_VDDO_res_M3_g N_VDDO_M3_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M1 U28_MPI2_drain N_U27_padr_M1_g N_VDDO_M1_s N_VDDO_M60_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M2 N_U28_MPI1_drain_M2_d N_U27_padr_M2_g U28_MPI2_drain N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M28 N_U15_U12_oenb_M28_d N_U15_U15_OUTSHIFT_M28_g N_VDDO_M28_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M28@2 N_U15_U12_oenb_M28@2_d N_U15_U15_OUTSHIFT_M28@2_g N_VDDO_M28_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M8 N_U15_pgate_M8_d N_U15_ISHF_M8_g N_VDDO_M8_s N_VDDO_M60_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M8@2 N_U15_pgate_M8@2_d N_U15_ISHF_M8@2_g N_VDDO_M8_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M29 N_U15_pgate_M8@2_d N_U15_U12_oenb_M29_g N_VDDO_M29_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M29@2 N_U15_pgate_M29@2_d N_U15_U12_oenb_M29@2_g N_VDDO_M29_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M9 N_U15_ngate_M9_d N_U15_U15_OUTSHIFT_M9_g N_U15_pgate_M9_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9@2 N_U15_ngate_M9_d N_U15_U15_OUTSHIFT_M9@2_g N_U15_pgate_M9@2_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M9@3 N_U15_ngate_M9@3_d N_U15_U15_OUTSHIFT_M9@3_g N_U15_pgate_M9@2_s
+ N_VDDO_M60_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M18 N_U15_U15_MPLL1_dr_M18_d N_U15_U15_OUTSHIFT_M18_g N_VDDO_M18_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M19 N_U15_U15_OUTSHIFT_M19_d N_U15_U15_MPLL1_dr_M19_g N_VDDO_M18_s N_VDDO_M60_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M10 N_U15_U14_MPLL1_dr_M10_d N_U15_ISHF_M10_g N_VDDO_M10_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U15_ISHF_M11_d N_U15_U14_MPLL1_dr_M11_g N_VDDO_M10_s N_VDDO_M60_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M16 N_U15_U14_MN1_drai_M16_d N_I_M16_g N_VDD_M16_s N_VDD_M16_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M16@2 N_U15_U14_MN1_drai_M16_d N_I_M16@2_g N_VDD_M16@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M24 N_U15_U15_MN1_drai_M24_d N_OEN_M24_g N_VDD_M16@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M24@2 N_U15_U15_MN1_drai_M24_d N_OEN_M24@2_g N_VDD_M24@2_s N_VDD_M16_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D17 N_VSS_M54_b N_I_D17_neg DN18  AREA=2.5e-13 PJ=2e-06
D25 N_VSS_M54_b N_OEN_D25_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM60 N_VSSO_RM60_pos N_net_m60_VSSO_res_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM3 N_net_m3_VDDO_res_RM3_pos N_VDDO_RM3_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM54 N_VDDO_RM54_pos N_net_m54_VDDO_res_RM54_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM59 N_VDDO_RM59_pos N_net_m59_VDDO_res_RM59_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_VSSO_RM4_pos N_net_m4_VSSO_res_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM55 N_net_m55_VSSO_res_RM55_pos N_VSSO_RM55_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U28_MPI2_drain 0 0.0289375f
*
.include "pc3t01.dist.sp.PC3T01.pxi"
*
.ends
*
*
* File: pc3t01u.dist.sp
* Created: Sun Jul  4 12:42:11 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t01u.dist.sp.pex"
.subckt pc3t01u  PAD I OEN VDD VSS VDDO VSSO 
* 
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M11 N_PAD_M12_d N_U27_U69$9_gate_M11_g N_VSSO_M11_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$9_gate_M12_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M14_d N_U27_U69$9_gate_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$9_gate_M14_g N_VSSO_M11_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$9_gate_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$9_gate_M16_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M17_d N_U15_ngate_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$9_gate_M17_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$9_gate_M18_g N_VSSO_M18_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U15_ngate_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U27_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M37_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$9_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M21 N_VDDO_M21_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M22 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M30_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M23_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M5 N_U27_padr_M5_d N_net_m5_VSSO_res_M5_g N_VSSO_M5_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5@2 N_U27_padr_M5@2_d N_net_m5_VSSO_res_M5@2_g N_VSSO_M5_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6 N_U29_MPI1_drain_M6_d N_U27_padr_M6_g N_VSSO_M6_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M4 N_U27_padr_M4_d N_net_m4_VDDO_res_M4_g N_VDDO_M4_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M2 U29_MPI2_drain N_U27_padr_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M3 N_U29_MPI1_drain_M3_d N_U27_padr_M3_g U29_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_net_m4_VDDO_res_RM4_pos N_VDDO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM5 N_VSSO_RM5_pos N_net_m5_VSSO_res_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_MPI2_drain 0 0.0289375f
*
.include "pc3t01u.dist.sp.PC3T01U.pxi"
*
.ends
*
*
* File: pc3t02d.dist.sp
* Created: Sun Jul  4 12:43:45 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t02d.dist.sp.pex"
.subckt pc3t02d  PAD I OEN VDD VSS VDDO VSSO 
* 
M67 N_U27_padr_M67_d N_net_m67_VDDO_res_M67_g U28_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M68 U28_U22_source N_net_m68_VDDO_res_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM67 N_net_m67_VDDO_res_RM67_pos N_VDDO_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM68 N_VDDO_RM67_neg N_net_m68_VDDO_res_RM68_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M65 N_U27_padr_M65_d N_net_m65_VSSO_res_M65_g N_VSSO_M65_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M65@2 N_U27_padr_M65@2_d N_net_m65_VSSO_res_M65@2_g N_VSSO_M65_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U29_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U29_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U29_MPI1_drain_M63_d N_U27_padr_M63_g U29_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM65 N_VSSO_RM65_pos N_net_m65_VSSO_res_RM65_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.361103f
c_2 U29_MPI2_drain 0 0.0169448f
*
.include "pc3t02d.dist.sp.PC3T02D.pxi"
*
.ends
*
*
* File: pc3t02.dist.sp
* Created: Sun Jul  4 12:43:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t02.dist.sp.pex"
.subckt pc3t02  PAD I OEN VDD VSS VDDO VSSO 
* 
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M65 N_U27_padr_M65_d N_net_m65_VSSO_res_M65_g N_VSSO_M65_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M65@2 N_U27_padr_M65@2_d N_net_m65_VSSO_res_M65@2_g N_VSSO_M65_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U28_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U28_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U28_MPI1_drain_M63_d N_U27_padr_M63_g U28_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM65 N_VSSO_RM65_pos N_net_m65_VSSO_res_RM65_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.361103f
c_2 U28_MPI2_drain 0 0.0169448f
*
.include "pc3t02.dist.sp.PC3T02.pxi"
*
.ends
*
*
* File: pc3t02u.dist.sp
* Created: Sun Jul  4 12:45:38 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t02u.dist.sp.pex"
.subckt pc3t02u  PAD I OEN VDD VSS VDDO VSSO 
* 
M11 N_PAD_M12_d N_U27_U69$7_gate_M11_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U27_U69$7_gate_M12_g N_VSSO_M12_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M13 N_PAD_M14_d N_U27_U69$7_gate_M13_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U27_U69$7_gate_M14_g N_VSSO_M11_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M16_d N_U27_U69$7_gate_M15_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U27_U69$7_gate_M16_g N_VSSO_M13_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M17_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U27_U69$7_gate_M17_g N_VSSO_M15_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M10_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M9_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M8_d N_U27_U69$7_gate_M18_g N_VSSO_M18_s N_VSSO_M12_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M12_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M67 N_U27_padr_M67_d N_net_m67_VSSO_res_M67_g N_VDDO_M67_s N_VDDO_M37_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U27_U72_pgate_M32_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U27_U72_pgate_M32@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U27_U72_pgate_M32@4_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR35 N_U27_U69$7_gate_R35_pos N_VSSO_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM67 N_net_m67_VSSO_res_RM67_pos N_VSSO_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U27_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M23 N_VDDO_M23_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M24 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M22_d N_U27_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_U27_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_U27_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U27_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U27_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U27_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U27_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U27_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M36 N_VDDO_M36_d N_net_m36_VDDO_res_M36_g N_U27_U71_UN_P_TOP_M36_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M65 N_U27_padr_M65_d N_net_m65_VSSO_res_M65_g N_VSSO_M65_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M65@2 N_U27_padr_M65@2_d N_net_m65_VSSO_res_M65@2_g N_VSSO_M65_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M66 N_U30_MPI1_drain_M66_d N_U27_padr_M66_g N_VSSO_M66_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M59 N_U15_U12_oenb_M59_d N_U15_U15_OUTSHIFT_M59_g N_VSSO_M59_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M38 N_U15_ngate_M38_d N_U15_ISHF_M38_g N_VSSO_M38_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_U15_ngate_M38_d N_U15_ISHF_M38@2_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M58 N_U15_ngate_M58_d N_U15_U15_OUTSHIFT_M58_g N_VSSO_M38@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M39 N_U15_pgate_M39_d N_U15_U12_oenb_M39_g N_U15_ngate_M39_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@2_g N_U15_ngate_M39_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M39@3 N_U15_pgate_M39@2_d N_U15_U12_oenb_M39@3_g N_U15_ngate_M39@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_OEN_M52_g N_VSSO_M52_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M54 N_VDDO_M54_d N_U15_U15_MN1_drai_M54_g N_U15_U15_MPLL1_dr_M54_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M52@2 N_U15_U15_MPLL1_dr_M52@2_d N_OEN_M52@2_g N_VSSO_M52_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MN1_drai_M53_g N_VSSO_M53_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M53@2 N_U15_U15_OUTSHIFT_M53@2_d N_U15_U15_MN1_drai_M53@2_g N_VSSO_M53_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M46 N_VDDO_M46_d N_U15_U14_MN1_drai_M46_g N_U15_U14_MPLL1_dr_M46_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M44 N_U15_U14_MPLL1_dr_M44_d N_I_M44_g N_VSSO_M44_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U15_U14_MPLL1_dr_M44@2_d N_I_M44@2_g N_VSSO_M44_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45 N_U15_ISHF_M45_d N_U15_U14_MN1_drai_M45_g N_VSSO_M45_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M45@2 N_U15_ISHF_M45@2_d N_U15_U14_MN1_drai_M45@2_g N_VSSO_M45_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U14_MN1_drai_M47_d N_I_M47_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M55 N_U15_U15_MN1_drai_M55_d N_OEN_M55_g N_VSS_M47_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M37 N_U27_U71_UN_P_TOP_M37_d N_net_m37_VSSO_res_M37_g N_VDDO_M37_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M37_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M37_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M37_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M64 N_U27_padr_M64_d N_net_m64_VDDO_res_M64_g N_VDDO_M64_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M62 U30_MPI2_drain N_U27_padr_M62_g N_VDDO_M62_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M63 N_U30_MPI1_drain_M63_d N_U27_padr_M63_g U30_MPI2_drain N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M60 N_U15_U12_oenb_M60_d N_U15_U15_OUTSHIFT_M60_g N_VDDO_M60_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60@2 N_U15_U12_oenb_M60@2_d N_U15_U15_OUTSHIFT_M60@2_g N_VDDO_M60_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U15_pgate_M40_d N_U15_ISHF_M40_g N_VDDO_M40_s N_VDDO_M37_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M40@2 N_U15_pgate_M40@2_d N_U15_ISHF_M40@2_g N_VDDO_M40_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M61 N_U15_pgate_M40@2_d N_U15_U12_oenb_M61_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M61@2 N_U15_pgate_M61@2_d N_U15_U12_oenb_M61@2_g N_VDDO_M61_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M41 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41_g N_U15_pgate_M41_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U15_ngate_M41_d N_U15_U15_OUTSHIFT_M41@2_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U15_ngate_M41@3_d N_U15_U15_OUTSHIFT_M41@3_g N_U15_pgate_M41@2_s
+ N_VDDO_M37_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M50 N_U15_U15_MPLL1_dr_M50_d N_U15_U15_OUTSHIFT_M50_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M51 N_U15_U15_OUTSHIFT_M51_d N_U15_U15_MPLL1_dr_M51_g N_VDDO_M50_s N_VDDO_M37_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MPLL1_dr_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M43 N_U15_ISHF_M43_d N_U15_U14_MPLL1_dr_M43_g N_VDDO_M42_s N_VDDO_M37_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M48 N_U15_U14_MN1_drai_M48_d N_I_M48_g N_VDD_M48_s N_VDD_M48_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M48@2 N_U15_U14_MN1_drai_M48_d N_I_M48@2_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56 N_U15_U15_MN1_drai_M56_d N_OEN_M56_g N_VDD_M48@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M56@2 N_U15_U15_MN1_drai_M56_d N_OEN_M56@2_g N_VDD_M56@2_s N_VDD_M48_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D49 N_VSS_M31_b N_I_D49_neg DN18  AREA=2.5e-13 PJ=2e-06
D57 N_VSS_M31_b N_OEN_D57_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM37 N_VSSO_RM37_pos N_net_m37_VSSO_res_RM37_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM64 N_net_m64_VDDO_res_RM64_pos N_VDDO_RM64_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM36 N_VDDO_RM36_pos N_net_m36_VDDO_res_RM36_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM65 N_VSSO_RM65_pos N_net_m65_VSSO_res_RM65_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.361103f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pc3t02u.dist.sp.PC3T02U.pxi"
*
.ends
*
*
* File: pc3t03d.dist.sp
* Created: Sun Jul  4 12:47:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t03d.dist.sp.pex"
.subckt pc3t03d  PAD I OEN VDD VSS VDDO VSSO 
* 
M69 N_U28_padr_M69_d N_net_m69_VDDO_res_M69_g U29_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U29_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pc3t03d.dist.sp.PC3T03D.pxi"
*
.ends
*
*
* File: pc3t03.dist.sp
* Created: Sun Jul  4 12:45:32 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t03.dist.sp.pex"
.subckt pc3t03  PAD I OEN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pc3t03.dist.sp.PC3T03.pxi"
*
.ends
*
*
* File: pc3t03u.dist.sp
* Created: Sun Jul  4 12:47:25 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t03u.dist.sp.pex"
.subckt pc3t03u  PAD I OEN VDD VSS VDDO VSSO 
* 
M37 N_PAD_M38_d N_U28_U42_r1_M37_g N_VSSO_M37_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M38_d N_U28_U42_r1_M38_g N_VSSO_M38_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M39 N_PAD_M40_d N_U28_U42_r1_M39_g N_VSSO_M39_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U28_U42_r1_M40_g N_VSSO_M37_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M41_d N_U15_ngate_M35_g N_VSSO_M35_s N_VSSO_M38_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M41_d N_U28_U42_r1_M41_g N_VSSO_M39_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M31 N_PAD_M36_d N_U17_ngate2_M31_g N_VSSO_M31_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U15_ngate_M36_g N_VSSO_M35_s N_VSSO_M38_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M32_d N_U28_ngate3_M33_g N_VSSO_M33_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_PAD_M32_d N_U17_ngate2_M32_g N_VSSO_M31_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M34_d N_U28_U42_r1_M42_g N_VSSO_M42_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M34_d N_U28_ngate3_M34_g N_VSSO_M33_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M63_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M56 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56_g N_U28_U72_pgate_M56_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M56@2 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56@2_g N_U28_U72_pgate_M56@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@3 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@3_g N_U28_U72_pgate_M56@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@4 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@4_g N_U28_U72_pgate_M56@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@5 N_U15_pgate_M56@5_d N_net_m56_VSSO_res_M56@5_g N_U28_U72_pgate_M56@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U28_U42_r1_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VSSO_res_RM69_pos N_VSSO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR57 N_noxref_2_R57_pos N_PAD_R57_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR58 N_noxref_2_R58_pos N_U28_padr_R58_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M49 N_VDDO_M49_d N_U28_U71_UN_P_TOP_M49_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M50 N_VDDO_M51_d N_U28_U71_UN_P_TOP_M50_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M48_d N_U28_U72_pgate_M43_g N_PAD_M43_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M44 N_VDDO_M44_d N_U28_U72_pgate_M44_g N_PAD_M43_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M51 N_VDDO_M51_d N_U28_U71_UN_P_TOP_M51_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U28_U71_UN_P_TOP_M52_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U28_U71_UN_P_TOP_M53_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U28_U71_UN_P_TOP_M54_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M45 N_VDDO_M54_d N_U28_U72_pgate_M45_g N_PAD_M45_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M46 N_VDDO_M46_d N_U28_U72_pgate_M46_g N_PAD_M45_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M47 N_VDDO_M46_d N_U28_U72_pgate_M47_g N_PAD_M47_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M48 N_VDDO_M48_d N_U28_U72_pgate_M48_g N_PAD_M47_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55_g N_U28_U72_pgate_M55_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M55@2 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55@2_g N_U28_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M55@3 N_U15_pgate_M55@3_d N_net_m55_VDDO_res_M55@3_g N_U28_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U28_U71_UN_P_TOP_M62_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M55_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M60 N_U28_ngate3_M60_d N_U17_ngatex_M60_g N_VSSO_M60_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M55_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M28 N_U15_U12_oenb_M28_d N_U15_U15_OUTSHIFT_M28_g N_VSSO_M28_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_U15_ngate_M7_d N_U15_ISHF_M7_g N_VSSO_M7_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M7@2 N_U15_ngate_M7_d N_U15_ISHF_M7@2_g N_VSSO_M7@2_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M27 N_U15_ngate_M27_d N_U15_U15_OUTSHIFT_M27_g N_VSSO_M7@2_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M8 N_U15_pgate_M8_d N_U15_U12_oenb_M8_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@2_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@3_g N_U15_ngate_M8@3_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M21 N_U15_U15_MPLL1_dr_M21_d N_OEN_M21_g N_VSSO_M21_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M23 N_VDDO_M23_d N_U15_U15_MN1_drai_M23_g N_U15_U15_MPLL1_dr_M23_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M21@2 N_U15_U15_MPLL1_dr_M21@2_d N_OEN_M21@2_g N_VSSO_M21_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22 N_U15_U15_OUTSHIFT_M22_d N_U15_U15_MN1_drai_M22_g N_VSSO_M22_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22@2 N_U15_U15_OUTSHIFT_M22@2_d N_U15_U15_MN1_drai_M22@2_g N_VSSO_M22_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M15 N_VDDO_M15_d N_U15_U14_MN1_drai_M15_g N_U15_U14_MPLL1_dr_M15_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U15_U14_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U15_U14_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U15_ISHF_M14_d N_U15_U14_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U15_ISHF_M14@2_d N_U15_U14_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U15_U14_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M24 N_U15_U15_MN1_drai_M24_d N_OEN_M24_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U28_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M63_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M63_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M59 N_U28_ngate3_M59_d N_U17_ngatex_M59_g N_U17_ngate2_M59_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M29 N_U15_U12_oenb_M29_d N_U15_U15_OUTSHIFT_M29_g N_VDDO_M29_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M29@2 N_U15_U12_oenb_M29@2_d N_U15_U15_OUTSHIFT_M29@2_g N_VDDO_M29_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M9 N_U15_pgate_M9_d N_U15_ISHF_M9_g N_VDDO_M9_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M9@2 N_U15_pgate_M9@2_d N_U15_ISHF_M9@2_g N_VDDO_M9_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M30 N_U15_pgate_M9@2_d N_U15_U12_oenb_M30_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M30@2 N_U15_pgate_M30@2_d N_U15_U12_oenb_M30@2_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M10 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10_g N_U15_pgate_M10_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M10@2 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10@2_g N_U15_pgate_M10@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M10@3 N_U15_ngate_M10@3_d N_U15_U15_OUTSHIFT_M10@3_g N_U15_pgate_M10@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M19 N_U15_U15_MPLL1_dr_M19_d N_U15_U15_OUTSHIFT_M19_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M20 N_U15_U15_OUTSHIFT_M20_d N_U15_U15_MPLL1_dr_M20_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U15_U14_MPLL1_dr_M11_d N_U15_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U15_ISHF_M12_d N_U15_U14_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M17 N_U15_U14_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U15_U14_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25 N_U15_U15_MN1_drai_M25_d N_OEN_M25_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25@2 N_U15_U15_MN1_drai_M25_d N_OEN_M25@2_g N_VDD_M25@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D18 N_VSS_M55_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
D26 N_VSS_M55_b N_OEN_D26_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM55 N_VDDO_RM55_pos N_net_m55_VDDO_res_RM55_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM56 N_net_m56_VSSO_res_RM56_pos N_VSSO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pc3t03u.dist.sp.PC3T03U.pxi"
*
.ends
*
*
* File: pc3t04d.dist.sp
* Created: Sun Jul  4 12:48:40 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t04d.dist.sp.pex"
.subckt pc3t04d  PAD I OEN VDD VSS VDDO VSSO 
* 
M69 N_U28_padr_M69_d N_net_m69_VDDO_res_M69_g U30_U22_source N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U30_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X36/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X36/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U31_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U31_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U31_MPI1_drain_M65_d N_U28_padr_M65_g U31_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U31_MPI2_drain 0 0.0169448f
*
.include "pc3t04d.dist.sp.PC3T04D.pxi"
*
.ends
*
*
* File: pc3t04.dist.sp
* Created: Sun Jul  4 12:48:33 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t04.dist.sp.pex"
.subckt pc3t04  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X32/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X32/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U29_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U29_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U29_MPI1_drain_M65_d N_U28_padr_M65_g U29_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U29_MPI2_drain 0 0.0169448f
*
.include "pc3t04.dist.sp.PC3T04.pxi"
*
.ends
*
*
* File: pc3t04u.dist.sp
* Created: Sun Jul  4 12:50:18 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t04u.dist.sp.pex"
.subckt pc3t04u  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M10_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M11_d N_U15_ngate_M9_g N_VSSO_M9_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M17_d N_U28_ngate3_M7_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M18_d N_U28_U42_r1_M16_g N_VSSO_M15_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M13_d N_U17_ngate2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M14_d N_U28_ngate3_M8_g N_VSSO_M7_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M20 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U28_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U15_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U28_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U15_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U15_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U28_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VSSO_res_RM69_pos N_VSSO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M10 N_PAD_M10_d N_U15_ngate_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U15_ngate_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U28_U42_r1_M18_g N_VSSO_M17_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U17_ngate2_M13_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U17_ngate2_M14_g N_VSSO_M13_s N_VSSO_M10_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_VDDO_M33_d N_U28_U71_UN_P_TOP_M33_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M34_g N_PAD_M33_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M32_d N_U28_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U28_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M35 N_VDDO_M35_d N_U28_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M36 N_VDDO_M36_d N_U28_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M36_d N_U28_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U28_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U28_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M35_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
XR21 N_X34/noxref_10_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_X34/noxref_10_R22_pos N_U28_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M19 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U28_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U15_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U15_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U28_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U28_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U28_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359779f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pc3t04u.dist.sp.PC3T04U.pxi"
*
.ends
*
*
* File: pc3t05d.dist.sp
* Created: Sun Jul  4 12:51:52 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t05d.dist.sp.pex"
.subckt pc3t05d  PAD I OEN VDD VSS VDDO VSSO 
* 
M69 N_U29_padr_M69_d N_net_m69_VDDO_res_M69_g U31_U22_source N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U31_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U32_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U32_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U32_MPI1_drain_M65_d N_U29_padr_M65_g U32_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U32_MPI2_drain 0 0.0169448f
*
.include "pc3t05d.dist.sp.PC3T05D.pxi"
*
.ends
*
*
* File: pc3t05.dist.sp
* Created: Sun Jul  4 12:50:12 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t05.dist.sp.pex"
.subckt pc3t05  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U31_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U31_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U31_MPI1_drain_M65_d N_U29_padr_M65_g U31_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U31_MPI2_drain 0 0.0169448f
*
.include "pc3t05.dist.sp.PC3T05.pxi"
*
.ends
*
*
* File: pc3t05u.dist.sp
* Created: Sun Jul  4 12:51:55 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3t05u.dist.sp.pex"
.subckt pc3t05u  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U32_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U32_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U32_MPI1_drain_M65_d N_U29_padr_M65_g U32_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U32_MPI2_drain 0 0.0169448f
*
.include "pc3t05u.dist.sp.PC3T05U.pxi"
*
.ends
*
*
* File: pc3x11.dist.sp
* Created: Sun Jul  4 12:53:42 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3x11.dist.sp.pex"
.subckt pc3x11  Z XIN EN XOUT VDD VSS VDDO VSSO 
* 
M94 N_U12_U19_source_M94_d N_U8_IN_M94_g N_VSS_M94_s N_VSS_M99_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M93 N_U12_U22_gate_M93_d N_U23_padr_M93_g N_U12_U19_source_M93_s N_VSS_M99_b
+ NHV L=3.6e-07 W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M35 N_XOUT_M33_d N_U23_U73$1_gate_M35_g N_VSSO_M38_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M36 N_XOUT_M34_d N_U23_U73$1_gate_M36_g N_VSSO_M43_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M2 N_U8_OUT_M2_d N_U8_IN_M2_g N_VSS_M2_s N_VSS_M99_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M4 N_U8_IN_M4_d N_EN_M4_g N_VSS_M2_s N_VSS_M99_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M91 N_U12_U22_drain_M91_d N_U12_U22_gate_M91_g N_VSS_M91_s N_VSS_M99_b N18
+ L=3.6e-07 W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M92 N_Z_M92_d N_U12_U22_drain_M92_g N_VSS_M92_s N_VSS_M99_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M92@2 N_Z_M92@2_d N_U12_U22_drain_M92@2_g N_VSS_M92_s N_VSS_M99_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M97 N_U12_U22_gate_M97_d N_U23_padr_M97_g N_VDD_M97_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M96 N_U12_U22_gate_M96_d N_U8_IN_M96_g N_VDD_M96_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M1 N_U8_OUT_M1_d N_U8_IN_M1_g N_VDD_M1_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M1@2 N_U8_OUT_M1_d N_U8_IN_M1@2_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.175e-05 AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3 N_U8_IN_M3_d N_EN_M3_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3@2 N_U8_IN_M3_d N_EN_M3@2_g N_VDD_M3@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M98 N_Z_M98_d N_U12_U22_drain_M98_g N_VDD_M98_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.4e-05 AD=8.68e-12 AS=6.1075e-12 PD=2.924e-05 PS=1.64675e-05
M98@2 N_Z_M98@2_d N_U12_U22_drain_M98@2_g N_VDD_M98_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.8e-05 AD=7.38e-12 AS=7.8525e-12 PD=1.882e-05 PS=2.11725e-05
M98@3 N_Z_M98@2_d N_U12_U22_drain_M98@3_g N_VDD_M98@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=7.38e-12 AS=7.38e-12 PD=1.882e-05 PS=1.882e-05
M95 N_U12_U22_drain_M95_d N_U12_U22_gate_M95_g N_VDD_M98@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=1.116e-11 AS=7.38e-12 PD=3.724e-05 PS=1.882e-05
D90 N_VSS_M99_b N_EN_D90_neg DN18  AREA=2.25e-12 PJ=6e-06
XR57 N_VDD_R57_pos N_U23_U37_r2_R57_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR55 N_VSS_R55_pos N_U23_U73$1_gate_R55_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M33 N_XOUT_M33_d N_U22_PADR_M33_g U23_MN4$1_drain N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M31 U23_MN4$1_drain N_U8_IN_M31_g N_VSSO_M31_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
M34 N_XOUT_M34_d N_U22_PADR_M34_g U23_MN4$0_drain N_VSSO_M33_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M32 U23_MN4$0_drain N_U8_IN_M32_g N_VSSO_M32_s N_VSSO_M33_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
XR72 N_VSS_R72_pos N_U22_U82_gate_R72_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR56 N_VDD_R56_pos U23_U72$1_gate RNWELLSTI2T w=2.1e-06 l=2.1e-06 
M37 N_XOUT_M37_d N_U23_U73$1_gate_M37_g N_VSSO_M37_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M38 N_XOUT_M37_d N_U23_U73$1_gate_M38_g N_VSSO_M38_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M39 N_XOUT_M39_d N_U23_U73$1_gate_M39_g N_VSSO_M39_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M40 N_XOUT_M39_d N_U23_U73$1_gate_M40_g N_VSSO_M37_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M41 N_XOUT_M41_d N_U23_U73$1_gate_M41_g N_VSSO_M41_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M42 N_XOUT_M41_d N_U23_U73$1_gate_M42_g N_VSSO_M39_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M43 N_XOUT_M43_d N_U23_U73$1_gate_M43_g N_VSSO_M43_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M44 N_XOUT_M43_d N_U23_U73$1_gate_M44_g N_VSSO_M41_s N_VSSO_M33_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M99 N_U23_padr_M99_d N_U12_U27$1_gate_M99_g N_VSS_M99_s N_VSS_M99_b N18 L=4e-07
+ W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
M100 N_U23_padr_M99_d N_U12_U27$1_gate_M100_g N_VSS_M100_s N_VSS_M99_b N18
+ L=4e-07 W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
XR53 N_U23_padr_R53_pos N_X0/X37/noxref_4_R53_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR54 N_X0/X37/noxref_4_R54_pos N_XOUT_R54_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M9 N_VDD_M9_d N_U23_U37_r2_M9_g U23_U82$9_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M19 U23_U82$9_source N_U23_U37_r2_M19_g N_XOUT_M19_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M20 U23_U82$8_source N_U23_U37_r2_M20_g N_XOUT_M19_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M10 N_VDD_M11_d N_U23_U37_r2_M10_g U23_U82$8_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M5 N_VDD_M18_d N_U8_OUT_M5_g U23_MP4$1_source N_VDD_M11_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M7 U23_MP4$1_source N_U22_PADR_M7_g N_XOUT_M7_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M8 U23_MP4$0_source N_U22_PADR_M8_g N_XOUT_M7_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M6 N_VDD_M6_d N_U8_OUT_M6_g U23_MP4$0_source N_VDD_M11_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M11 N_VDD_M11_d N_U23_U37_r2_M11_g U23_U82$7_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M21 U23_U82$7_source N_U23_U37_r2_M21_g N_XOUT_M21_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M22 U23_U82$6_source N_U23_U37_r2_M22_g N_XOUT_M21_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M12 N_VDD_M12_d N_U23_U37_r2_M12_g U23_U82$6_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M13 N_VDD_M12_d N_U23_U37_r2_M13_g U23_U82$5_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M23 U23_U82$5_source N_U23_U37_r2_M23_g N_XOUT_M23_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M24 U23_U82$4_source N_U23_U37_r2_M24_g N_XOUT_M23_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M14 N_VDD_M14_d N_U23_U37_r2_M14_g U23_U82$4_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M15 N_VDD_M14_d N_U23_U37_r2_M15_g U23_U82$3_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M25 U23_U82$3_source N_U23_U37_r2_M25_g N_XOUT_M25_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M26 U23_U82$2_source N_U23_U37_r2_M26_g N_XOUT_M25_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M16 N_VDD_M16_d N_U23_U37_r2_M16_g U23_U82$2_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M17 N_VDD_M16_d N_U23_U37_r2_M17_g U23_U82$1_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M27 U23_U82$1_source N_U23_U37_r2_M27_g N_XOUT_M27_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M28 U23_U82$0_source N_U23_U37_r2_M28_g N_XOUT_M27_s N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M18 N_VDD_M18_d N_U23_U37_r2_M18_g U23_U82$0_source N_VDD_M11_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M76 N_XIN_M82_d N_U22_R_PULLDONW_r_M76_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M77 N_XIN_M83_d N_U22_R_PULLDONW_r_M77_g N_VSSO_M77_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M78 N_XIN_M84_d N_U22_R_PULLDONW_r_M78_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M79 N_XIN_M85_d N_U22_R_PULLDONW_r_M79_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M80 N_XIN_M86_d N_U22_R_PULLDONW_r_M80_g N_VSSO_M80_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M81 N_XIN_M87_d N_U22_R_PULLDONW_r_M81_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
MPCL N_U22_PADR_MPCL_d N_RU1_MPCL_g N_VDD_MPCL_s N_VDD_M1_b P18 L=5e-07 W=2e-05
+ AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
MPCL@2 N_U22_PADR_MPCL_d N_RU1_MPCL@2_g N_VDD_MPCL@2_s N_VDD_M1_b P18 L=5e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
D89@2 N_VSS_D89@2_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@3 N_VSS_D89@3_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@4 N_VSS_D89@4_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@5 N_VSS_D89@5_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@6 N_VSS_D89@6_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@7 N_VSS_D89@7_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89 N_VSS_D89_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@2 N_VSSO_D88@2_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@3 N_VSSO_D88@3_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@4 N_VSSO_D88@4_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@5 N_VSSO_D88@5_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@6 N_VSSO_D88@6_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@7 N_VSSO_D88@7_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88 N_VSSO_D88_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XRPUP1 N_RU1_RPUP1_pos N_VDD_RPUP1_neg RPMPOLY2T w=2e-06 l=8e-06 
XR73 N_U22_R_PULLDONW_r_R73_pos N_VSSO_R73_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06
+ 
XR74 N_U22_U79$3_gate_R74_pos N_VDDO_R74_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR102 N_VSS_R102_pos N_U12_U27$1_gate_R102_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR70 N_U22_PADR_R70_pos N_X1/X29/noxref_4_R70_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR71 N_X1/X29/noxref_4_R71_pos N_XIN_R71_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M82 N_XIN_M82_d N_U22_R_PULLDONW_r_M82_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M83 N_XIN_M83_d N_U22_R_PULLDONW_r_M83_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M84 N_XIN_M84_d N_U22_R_PULLDONW_r_M84_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M85 N_XIN_M85_d N_U22_R_PULLDONW_r_M85_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M86 N_XIN_M86_d N_U22_R_PULLDONW_r_M86_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M87 N_XIN_M87_d N_U22_R_PULLDONW_r_M87_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M75 N_U22_PADR_M75_d N_U22_U82_gate_M75_g N_VSS_M75_s N_VSS_M75_b N18 L=4e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M75@2 N_U22_PADR_M75_d N_U22_U82_gate_M75@2_g N_VSS_M75@2_s N_VSS_M75_b N18
+ L=4e-07 W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M58 N_VDDO_M58_d N_U22_U79$3_gate_M58_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M59 N_VDDO_M62_d N_U22_U79$3_gate_M59_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M60 N_VDDO_M69_d N_U22_U79$3_gate_M60_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M61 N_VDDO_M61_d N_U22_U79$3_gate_M61_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M62 N_VDDO_M62_d N_U22_U79$3_gate_M62_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M63 N_VDDO_M63_d N_U22_U79$3_gate_M63_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M64 N_VDDO_M63_d N_U22_U79$3_gate_M64_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M65 N_VDDO_M65_d N_U22_U79$3_gate_M65_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M66 N_VDDO_M65_d N_U22_U79$3_gate_M66_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M67 N_VDDO_M67_d N_U22_U79$3_gate_M67_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M68 N_VDDO_M67_d N_U22_U79$3_gate_M68_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M69 N_VDDO_M69_d N_U22_U79$3_gate_M69_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U23_U72$1_gate 0 39.4256f
c_2 U23_MN4$1_drain 0 0.0877515f
c_3 U23_MN4$0_drain 0 0.0877515f
c_4 U23_U82$9_source 0 0.01206f
c_5 U23_U82$8_source 0 0.01206f
c_6 U23_MP4$1_source 0 0.0268754f
c_7 U23_MP4$0_source 0 0.0270855f
c_8 U23_U82$7_source 0 0.0116103f
c_9 U23_U82$6_source 0 0.0116103f
c_10 U23_U82$5_source 0 0.0116103f
c_11 U23_U82$4_source 0 0.0116103f
c_12 U23_U82$3_source 0 0.0116103f
c_13 U23_U82$2_source 0 0.0116103f
c_14 U23_U82$1_source 0 0.0116103f
c_15 U23_U82$0_source 0 0.0116103f
*
.include "pc3x11.dist.sp.PC3X11.pxi"
*
.ends
*
*
* File: pc3x12.dist.sp
* Created: Sun Jul  4 12:53:32 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3x12.dist.sp.pex"
.subckt pc3x12  Z XIN EN XOUT VDD VSS VDDO VSSO 
* 
M93 N_U12_U19_source_M93_d N_U8_IN_M93_g N_VSS_M93_s N_VSS_M98_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M92 N_U12_U22_gate_M92_d N_U23_padr_M92_g N_U12_U19_source_M92_s N_VSS_M98_b
+ NHV L=3.6e-07 W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M2 N_U8_OUT_M2_d N_U8_IN_M2_g N_VSS_M2_s N_VSS_M98_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M4 N_U8_IN_M4_d N_EN_M4_g N_VSS_M2_s N_VSS_M98_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M90 N_U12_U22_drain_M90_d N_U12_U22_gate_M90_g N_VSS_M90_s N_VSS_M98_b N18
+ L=3.6e-07 W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M91 N_Z_M91_d N_U12_U22_drain_M91_g N_VSS_M91_s N_VSS_M98_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M91@2 N_Z_M91@2_d N_U12_U22_drain_M91@2_g N_VSS_M91_s N_VSS_M98_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M96 N_U12_U22_gate_M96_d N_U23_padr_M96_g N_VDD_M96_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M95 N_U12_U22_gate_M95_d N_U8_IN_M95_g N_VDD_M95_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M1 N_U8_OUT_M1_d N_U8_IN_M1_g N_VDD_M1_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M1@2 N_U8_OUT_M1_d N_U8_IN_M1@2_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.175e-05 AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3 N_U8_IN_M3_d N_EN_M3_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3@2 N_U8_IN_M3_d N_EN_M3@2_g N_VDD_M3@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M97 N_Z_M97_d N_U12_U22_drain_M97_g N_VDD_M97_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.4e-05 AD=8.68e-12 AS=6.1075e-12 PD=2.924e-05 PS=1.64675e-05
M97@2 N_Z_M97@2_d N_U12_U22_drain_M97@2_g N_VDD_M97_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.8e-05 AD=7.38e-12 AS=7.8525e-12 PD=1.882e-05 PS=2.11725e-05
M97@3 N_Z_M97@2_d N_U12_U22_drain_M97@3_g N_VDD_M97@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=7.38e-12 AS=7.38e-12 PD=1.882e-05 PS=1.882e-05
M94 N_U12_U22_drain_M94_d N_U12_U22_gate_M94_g N_VDD_M97@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=1.116e-11 AS=7.38e-12 PD=3.724e-05 PS=1.882e-05
D102 N_VSS_M98_b N_EN_D102_neg DN18  AREA=2.25e-12 PJ=6e-06
M37 N_XOUT_M37_d N_U22_PADR_M37_g U23_MN4$3_drain N_VSSO_M41_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M33 U23_MN4$3_drain N_U8_IN_M33_g N_VSSO_M33_s N_VSSO_M41_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
M38 N_XOUT_M32_d N_U22_PADR_M38_g U23_MN4$2_drain N_VSSO_M41_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M34 U23_MN4$2_drain N_U8_IN_M34_g N_VSSO_M34_s N_VSSO_M41_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M39 N_XOUT_M39_d N_U22_PADR_M39_g U23_MN4$1_drain N_VSSO_M41_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M35 U23_MN4$1_drain N_U8_IN_M35_g N_VSSO_M34_s N_VSSO_M41_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M40 N_XOUT_M39_d N_U22_PADR_M40_g U23_MN4$0_drain N_VSSO_M41_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M36 U23_MN4$0_drain N_U8_IN_M36_g N_VSSO_M36_s N_VSSO_M41_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
M31 N_XOUT_M37_d N_U23_U73$1_gate_M31_g N_VSSO_M42_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M32 N_XOUT_M32_d N_U23_U73$1_gate_M32_g N_VSSO_M45_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M41 N_XOUT_M41_d N_U23_U73$1_gate_M41_g N_VSSO_M41_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M42 N_XOUT_M41_d N_U23_U73$1_gate_M42_g N_VSSO_M42_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M43 N_XOUT_M43_d N_U23_U73$1_gate_M43_g N_VSSO_M43_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M44 N_XOUT_M43_d N_U23_U73$1_gate_M44_g N_VSSO_M41_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M45 N_XOUT_M45_d N_U23_U73$1_gate_M45_g N_VSSO_M45_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M46 N_XOUT_M45_d N_U23_U73$1_gate_M46_g N_VSSO_M43_s N_VSSO_M41_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDD_M15_d N_U23_U37_r2_M15_g U23_U82$6_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M22 U23_U82$6_source N_U23_U37_r2_M22_g N_XOUT_M22_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M23 U23_U82$5_source N_U23_U37_r2_M23_g N_XOUT_M22_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M16 N_VDD_M17_d N_U23_U37_r2_M16_g U23_U82$5_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M5 N_VDD_M9_d N_U8_OUT_M5_g U23_MP4$4_source N_VDD_M17_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M10 U23_MP4$4_source N_U22_PADR_M10_g N_XOUT_M10_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M11 U23_MP4$3_source N_U22_PADR_M11_g N_XOUT_M10_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M6 N_VDD_M6_d N_U8_OUT_M6_g U23_MP4$3_source N_VDD_M17_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M17 N_VDD_M17_d N_U23_U37_r2_M17_g U23_U82$4_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M24 U23_U82$4_source N_U23_U37_r2_M24_g N_XOUT_M24_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M25 U23_U82$3_source N_U23_U37_r2_M25_g N_XOUT_M24_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M18 N_VDD_M18_d N_U23_U37_r2_M18_g U23_U82$3_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M19 N_VDD_M18_d N_U23_U37_r2_M19_g U23_U82$2_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M26 U23_U82$2_source N_U23_U37_r2_M26_g N_XOUT_M26_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M27 U23_U82$1_source N_U23_U37_r2_M27_g N_XOUT_M26_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M20 N_VDD_M20_d N_U23_U37_r2_M20_g U23_U82$1_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M21 N_VDD_M20_d N_U23_U37_r2_M21_g U23_U82$0_source N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M28 U23_U82$0_source N_U23_U37_r2_M28_g N_XOUT_M28_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M12 U23_MP4$2_source N_U22_PADR_M12_g N_XOUT_M28_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M7 N_VDD_M7_d N_U8_OUT_M7_g U23_MP4$2_source N_VDD_M17_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M8 N_VDD_M7_d N_U8_OUT_M8_g U23_MP4$1_source N_VDD_M17_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M13 U23_MP4$1_source N_U22_PADR_M13_g N_XOUT_M13_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M14 U23_MP4$0_source N_U22_PADR_M14_g N_XOUT_M13_s N_VDD_M17_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M9 N_VDD_M9_d N_U8_OUT_M9_g U23_MP4$0_source N_VDD_M17_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
XR53 N_U23_padr_R53_pos N_X0/X22/noxref_4_R53_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR54 N_X0/X22/noxref_4_R54_pos N_XOUT_R54_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M98 N_U23_padr_M98_d N_U12_U27$1_gate_M98_g N_VSS_M98_s N_VSS_M98_b N18 L=4e-07
+ W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
M99 N_U23_padr_M98_d N_U12_U27$1_gate_M99_g N_VSS_M99_s N_VSS_M98_b N18 L=4e-07
+ W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
XR72 N_VSS_R72_pos N_U22_U82_gate_R72_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR56 N_VDD_R56_pos U23_U72$1_gate RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR57 N_VDD_R57_pos N_U23_U37_r2_R57_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR55 N_VSS_R55_pos N_U23_U73$1_gate_R55_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M76 N_XIN_M82_d N_U22_R_PULLDONW_r_M76_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M77 N_XIN_M83_d N_U22_R_PULLDONW_r_M77_g N_VSSO_M77_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M78 N_XIN_M84_d N_U22_R_PULLDONW_r_M78_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M79 N_XIN_M85_d N_U22_R_PULLDONW_r_M79_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M80 N_XIN_M86_d N_U22_R_PULLDONW_r_M80_g N_VSSO_M80_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M81 N_XIN_M87_d N_U22_R_PULLDONW_r_M81_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
MPCL N_U22_PADR_MPCL_d N_RU1_MPCL_g N_VDD_MPCL_s N_VDD_M1_b P18 L=5e-07 W=2e-05
+ AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
MPCL@2 N_U22_PADR_MPCL_d N_RU1_MPCL@2_g N_VDD_MPCL@2_s N_VDD_M1_b P18 L=5e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
D89@2 N_VSS_D89@2_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@3 N_VSS_D89@3_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@4 N_VSS_D89@4_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@5 N_VSS_D89@5_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@6 N_VSS_D89@6_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@7 N_VSS_D89@7_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89 N_VSS_D89_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@2 N_VSSO_D88@2_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@3 N_VSSO_D88@3_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@4 N_VSSO_D88@4_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@5 N_VSSO_D88@5_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@6 N_VSSO_D88@6_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@7 N_VSSO_D88@7_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88 N_VSSO_D88_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XRPUP1 N_RU1_RPUP1_pos N_VDD_RPUP1_neg RPMPOLY2T w=2e-06 l=8e-06 
XR70 N_U22_PADR_R70_pos N_X1/X25/noxref_4_R70_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR71 N_X1/X25/noxref_4_R71_pos N_XIN_R71_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR101 N_VSS_R101_pos N_U12_U27$1_gate_R101_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR73 N_U22_R_PULLDONW_r_R73_pos N_VSSO_R73_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06
+ 
XR74 N_U22_U79$3_gate_R74_pos N_VDDO_R74_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M82 N_XIN_M82_d N_U22_R_PULLDONW_r_M82_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M83 N_XIN_M83_d N_U22_R_PULLDONW_r_M83_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M84 N_XIN_M84_d N_U22_R_PULLDONW_r_M84_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M85 N_XIN_M85_d N_U22_R_PULLDONW_r_M85_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M86 N_XIN_M86_d N_U22_R_PULLDONW_r_M86_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M87 N_XIN_M87_d N_U22_R_PULLDONW_r_M87_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M75 N_U22_PADR_M75_d N_U22_U82_gate_M75_g N_VSS_M75_s N_VSS_M75_b N18 L=4e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M75@2 N_U22_PADR_M75_d N_U22_U82_gate_M75@2_g N_VSS_M75@2_s N_VSS_M75_b N18
+ L=4e-07 W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M58 N_VDDO_M58_d N_U22_U79$3_gate_M58_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M59 N_VDDO_M62_d N_U22_U79$3_gate_M59_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M60 N_VDDO_M69_d N_U22_U79$3_gate_M60_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M61 N_VDDO_M61_d N_U22_U79$3_gate_M61_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M62 N_VDDO_M62_d N_U22_U79$3_gate_M62_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M63 N_VDDO_M63_d N_U22_U79$3_gate_M63_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M64 N_VDDO_M63_d N_U22_U79$3_gate_M64_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M65 N_VDDO_M65_d N_U22_U79$3_gate_M65_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M66 N_VDDO_M65_d N_U22_U79$3_gate_M66_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M67 N_VDDO_M67_d N_U22_U79$3_gate_M67_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M68 N_VDDO_M67_d N_U22_U79$3_gate_M68_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M69 N_VDDO_M69_d N_U22_U79$3_gate_M69_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U23_U72$1_gate 0 37.5792f
c_2 U23_MN4$3_drain 0 0.0877515f
c_3 U23_MN4$2_drain 0 0.0877559f
c_4 U23_MN4$1_drain 0 0.0877559f
c_5 U23_MN4$0_drain 0 0.088001f
c_6 U23_U82$6_source 0 0.01206f
c_7 U23_U82$5_source 0 0.01206f
c_8 U23_MP4$4_source 0 0.0269009f
c_9 U23_MP4$3_source 0 0.0270855f
c_10 U23_U82$4_source 0 0.0116103f
c_11 U23_U82$3_source 0 0.0116103f
c_12 U23_U82$2_source 0 0.0116103f
c_13 U23_U82$1_source 0 0.0116103f
c_14 U23_U82$0_source 0 0.0116103f
c_15 U23_MP4$2_source 0 0.0269009f
c_16 U23_MP4$1_source 0 0.0269009f
c_17 U23_MP4$0_source 0 0.0269009f
*
.include "pc3x12.dist.sp.PC3X12.pxi"
*
.ends
*
*
* File: pc3x13.dist.sp
* Created: Sun Jul  4 12:55:13 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pc3x13.dist.sp.pex"
.subckt pc3x13  Z XIN EN XOUT VDD VSS VDDO VSSO 
* 
M94 N_U12_U19_source_M94_d N_U8_IN_M94_g N_VSS_M94_s N_VSS_M99_b NHV L=3.6e-07
+ W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M93 N_U12_U22_gate_M93_d N_U23_padr_M93_g N_U12_U19_source_M93_s N_VSS_M99_b
+ NHV L=3.6e-07 W=4e-06 AD=2.48e-12 AS=2.48e-12 PD=9.24e-06 PS=9.24e-06
M2 N_U8_OUT_M2_d N_U8_IN_M2_g N_VSS_M2_s N_VSS_M99_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M4 N_U8_IN_M4_d N_EN_M4_g N_VSS_M2_s N_VSS_M99_b N18 L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M91 N_U12_U22_drain_M91_d N_U12_U22_gate_M91_g N_VSS_M91_s N_VSS_M99_b N18
+ L=3.6e-07 W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M92 N_Z_M92_d N_U12_U22_drain_M92_g N_VSS_M92_s N_VSS_M99_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M92@2 N_Z_M92@2_d N_U12_U22_drain_M92@2_g N_VSS_M92_s N_VSS_M99_b N18 L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M97 N_U12_U22_gate_M97_d N_U23_padr_M97_g N_VDD_M97_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M96 N_U12_U22_gate_M96_d N_U8_IN_M96_g N_VDD_M96_s N_VDD_M1_b PHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M1 N_U8_OUT_M1_d N_U8_IN_M1_g N_VDD_M1_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M1@2 N_U8_OUT_M1_d N_U8_IN_M1@2_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.175e-05 AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3 N_U8_IN_M3_d N_EN_M3_g N_VDD_M1@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=4.8175e-12 PD=1.257e-05 PS=1.257e-05
M3@2 N_U8_IN_M3_d N_EN_M3@2_g N_VDD_M3@2_s N_VDD_M1_b P18 L=3.6e-07 W=1.175e-05
+ AD=4.8175e-12 AS=7.285e-12 PD=1.257e-05 PS=2.474e-05
M98 N_Z_M98_d N_U12_U22_drain_M98_g N_VDD_M98_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.4e-05 AD=8.68e-12 AS=6.1075e-12 PD=2.924e-05 PS=1.64675e-05
M98@2 N_Z_M98@2_d N_U12_U22_drain_M98@2_g N_VDD_M98_s N_VDD_M1_b P18 L=3.6e-07
+ W=1.8e-05 AD=7.38e-12 AS=7.8525e-12 PD=1.882e-05 PS=2.11725e-05
M98@3 N_Z_M98@2_d N_U12_U22_drain_M98@3_g N_VDD_M98@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=7.38e-12 AS=7.38e-12 PD=1.882e-05 PS=1.882e-05
M95 N_U12_U22_drain_M95_d N_U12_U22_gate_M95_g N_VDD_M98@3_s N_VDD_M1_b P18
+ L=3.6e-07 W=1.8e-05 AD=1.116e-11 AS=7.38e-12 PD=3.724e-05 PS=1.882e-05
D90 N_VSS_M99_b N_EN_D90_neg DN18  AREA=2.25e-12 PJ=6e-06
M39 N_XOUT_M39_d N_U22_PADR_M39_g U23_MN4$5_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M33 U23_MN4$5_drain N_U8_IN_M33_g N_VSSO_M33_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
M40 N_XOUT_M32_d N_U22_PADR_M40_g U23_MN4$4_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=8.97e-11 AS=6.6e-12 PD=3.598e-05 PS=3.044e-05
M34 U23_MN4$4_drain N_U8_IN_M34_g N_VSSO_M34_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M41 N_XOUT_M41_d N_U22_PADR_M41_g U23_MN4$3_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M35 U23_MN4$3_drain N_U8_IN_M35_g N_VSSO_M34_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M42 N_XOUT_M41_d N_U22_PADR_M42_g U23_MN4$2_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M36 U23_MN4$2_drain N_U8_IN_M36_g N_VSSO_M36_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M43 N_XOUT_M43_d N_U22_PADR_M43_g U23_MN4$1_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M37 U23_MN4$1_drain N_U8_IN_M37_g N_VSSO_M36_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=2.28e-11 PD=3.044e-05 PS=3.152e-05
M44 N_XOUT_M43_d N_U22_PADR_M44_g U23_MN4$0_drain N_VSSO_M45_b NHV L=5e-07
+ W=3e-05 AD=7.56e-11 AS=6.6e-12 PD=3.504e-05 PS=3.044e-05
M38 U23_MN4$0_drain N_U8_IN_M38_g N_VSSO_M38_s N_VSSO_M45_b NHV L=5e-07 W=3e-05
+ AD=6.6e-12 AS=3.81e-11 PD=3.044e-05 PS=6.254e-05
M31 N_XOUT_M39_d N_U23_U73$1_gate_M31_g N_VSSO_M46_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M32 N_XOUT_M32_d N_U23_U73$1_gate_M32_g N_VSSO_M47_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=8.97e-11 AS=2.58e-11 PD=3.598e-05 PS=3.172e-05
M45 N_XOUT_M45_d N_U23_U73$1_gate_M45_g N_VSSO_M45_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M46 N_XOUT_M45_d N_U23_U73$1_gate_M46_g N_VSSO_M46_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M47 N_XOUT_M47_d N_U23_U73$1_gate_M47_g N_VSSO_M47_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M48 N_XOUT_M47_d N_U23_U73$1_gate_M48_g N_VSSO_M45_s N_VSSO_M45_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M21 N_VDD_M21_d N_U23_U37_r2_M21_g U23_U85$3_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M25 U23_U85$3_source N_U23_U37_r2_M25_g N_XOUT_M25_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M26 U23_U85$2_source N_U23_U37_r2_M26_g N_XOUT_M25_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M22 N_VDD_M22_d N_U23_U37_r2_M22_g U23_U85$2_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M23 N_VDD_M22_d N_U23_U37_r2_M23_g U23_U85$1_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M27 U23_U85$1_source N_U23_U37_r2_M27_g N_XOUT_M27_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M28 U23_U85$0_source N_U23_U37_r2_M28_g N_XOUT_M27_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M24 N_VDD_M7_d N_U23_U37_r2_M24_g U23_U85$0_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M5 N_VDD_M12_d N_U8_OUT_M5_g U23_MP4$7_source N_VDD_M7_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M13 U23_MP4$7_source N_U22_PADR_M13_g N_XOUT_M13_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M14 U23_MP4$6_source N_U22_PADR_M14_g N_XOUT_M13_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M6 N_VDD_M6_d N_U8_OUT_M6_g U23_MP4$6_source N_VDD_M7_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.04e-11 PD=0.00010684 PS=5.24e-05
M7 N_VDD_M7_d N_U8_OUT_M7_g U23_MP4$5_source N_VDD_M7_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M15 U23_MP4$5_source N_U22_PADR_M15_g N_XOUT_M15_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M16 U23_MP4$4_source N_U22_PADR_M16_g N_XOUT_M15_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M8 N_VDD_M8_d N_U8_OUT_M8_g U23_MP4$4_source N_VDD_M7_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M9 N_VDD_M8_d N_U8_OUT_M9_g U23_MP4$3_source N_VDD_M7_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M17 U23_MP4$3_source N_U22_PADR_M17_g N_XOUT_M17_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M18 U23_MP4$2_source N_U22_PADR_M18_g N_XOUT_M17_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M10 N_VDD_M10_d N_U8_OUT_M10_g U23_MP4$2_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M11 N_VDD_M10_d N_U8_OUT_M11_g U23_MP4$1_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
M19 U23_MP4$1_source N_U22_PADR_M19_g N_XOUT_M19_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M20 U23_MP4$0_source N_U22_PADR_M20_g N_XOUT_M19_s N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=1.04e-11 AS=1.2064e-10 PD=5.24e-05 PS=5.664e-05
M12 N_VDD_M12_d N_U8_OUT_M12_g U23_MP4$0_source N_VDD_M7_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.04e-11 PD=5.382e-05 PS=5.24e-05
XR53 N_U23_padr_R53_pos N_X0/X22/noxref_4_R53_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR54 N_X0/X22/noxref_4_R54_pos N_XOUT_R54_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M99 N_U23_padr_M99_d N_U12_U27$1_gate_M99_g N_VSS_M99_s N_VSS_M99_b N18 L=4e-07
+ W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
M100 N_U23_padr_M99_d N_U12_U27$1_gate_M100_g N_VSS_M100_s N_VSS_M99_b N18
+ L=4e-07 W=1.5e-05 AD=5.04e-11 AS=2.145e-11 PD=2.172e-05 PS=3.286e-05
XR72 N_VSS_R72_pos N_U22_U82_gate_R72_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR56 N_VDD_R56_pos U23_U72$1_gate RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR57 N_VDD_R57_pos N_U23_U37_r2_R57_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR55 N_VSS_R55_pos N_U23_U73$1_gate_R55_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M76 N_XIN_M82_d N_U22_R_PULLDONW_r_M76_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M77 N_XIN_M83_d N_U22_R_PULLDONW_r_M77_g N_VSSO_M77_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M78 N_XIN_M84_d N_U22_R_PULLDONW_r_M78_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M79 N_XIN_M85_d N_U22_R_PULLDONW_r_M79_g N_VSSO_M76_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M80 N_XIN_M86_d N_U22_R_PULLDONW_r_M80_g N_VSSO_M80_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M81 N_XIN_M87_d N_U22_R_PULLDONW_r_M81_g N_VSSO_M78_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
MPCL N_U22_PADR_MPCL_d N_RU1_MPCL_g N_VDD_MPCL_s N_VDD_M1_b P18 L=5e-07 W=2e-05
+ AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
MPCL@2 N_U22_PADR_MPCL_d N_RU1_MPCL@2_g N_VDD_MPCL@2_s N_VDD_M1_b P18 L=5e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
D89@2 N_VSS_D89@2_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@3 N_VSS_D89@3_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@4 N_VSS_D89@4_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@5 N_VSS_D89@5_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@6 N_VSS_D89@6_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89@7 N_VSS_D89@7_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D89 N_VSS_D89_pos N_VSSO_D89@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@2 N_VSSO_D88@2_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@3 N_VSSO_D88@3_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@4 N_VSSO_D88@4_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@5 N_VSSO_D88@5_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@6 N_VSSO_D88@6_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88@7 N_VSSO_D88@7_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D88 N_VSSO_D88_pos N_VSS_D88@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XRPUP1 N_RU1_RPUP1_pos N_VDD_RPUP1_neg RPMPOLY2T w=2e-06 l=8e-06 
XR70 N_U22_PADR_R70_pos N_X1/X25/noxref_4_R70_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR71 N_X1/X25/noxref_4_R71_pos N_XIN_R71_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR102 N_VSS_R102_pos N_U12_U27$1_gate_R102_neg RNWELLSTI2T w=2.1e-06 l=2.1e-06 
XR73 N_U22_R_PULLDONW_r_R73_pos N_VSSO_R73_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06
+ 
XR74 N_U22_U79$3_gate_R74_pos N_VDDO_R74_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M82 N_XIN_M82_d N_U22_R_PULLDONW_r_M82_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M83 N_XIN_M83_d N_U22_R_PULLDONW_r_M83_g N_VSSO_M82_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M84 N_XIN_M84_d N_U22_R_PULLDONW_r_M84_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M85 N_XIN_M85_d N_U22_R_PULLDONW_r_M85_g N_VSSO_M84_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M86 N_XIN_M86_d N_U22_R_PULLDONW_r_M86_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M87 N_XIN_M87_d N_U22_R_PULLDONW_r_M87_g N_VSSO_M86_s N_VSSO_M82_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M75 N_U22_PADR_M75_d N_U22_U82_gate_M75_g N_VSS_M75_s N_VSS_M75_b N18 L=4e-07
+ W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M75@2 N_U22_PADR_M75_d N_U22_U82_gate_M75@2_g N_VSS_M75@2_s N_VSS_M75_b N18
+ L=4e-07 W=2e-05 AD=4.66e-11 AS=4.97e-11 PD=2.466e-05 PS=4.497e-05
M58 N_VDDO_M58_d N_U22_U79$3_gate_M58_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M59 N_VDDO_M62_d N_U22_U79$3_gate_M59_g N_XIN_M58_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M60 N_VDDO_M69_d N_U22_U79$3_gate_M60_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M61 N_VDDO_M61_d N_U22_U79$3_gate_M61_g N_XIN_M60_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M62 N_VDDO_M62_d N_U22_U79$3_gate_M62_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M63 N_VDDO_M63_d N_U22_U79$3_gate_M63_g N_XIN_M62_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M64 N_VDDO_M63_d N_U22_U79$3_gate_M64_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M65 N_VDDO_M65_d N_U22_U79$3_gate_M65_g N_XIN_M64_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M66 N_VDDO_M65_d N_U22_U79$3_gate_M66_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M67 N_VDDO_M67_d N_U22_U79$3_gate_M67_g N_XIN_M66_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M68 N_VDDO_M67_d N_U22_U79$3_gate_M68_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M69 N_VDDO_M69_d N_U22_U79$3_gate_M69_g N_XIN_M68_s N_VDDO_M62_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U23_U72$1_gate 0 35.4454f
c_2 U23_MN4$5_drain 0 0.0877515f
c_3 U23_MN4$4_drain 0 0.0877559f
c_4 U23_MN4$3_drain 0 0.0877559f
c_5 U23_MN4$2_drain 0 0.0877559f
c_6 U23_MN4$1_drain 0 0.0877559f
c_7 U23_MN4$0_drain 0 0.088001f
c_8 U23_U85$3_source 0 0.01206f
c_9 U23_U85$2_source 0 0.01206f
c_10 U23_U85$1_source 0 0.0116103f
c_11 U23_U85$0_source 0 0.0116103f
c_12 U23_MP4$7_source 0 0.0268771f
c_13 U23_MP4$6_source 0 0.0270855f
c_14 U23_MP4$5_source 0 0.0268771f
c_15 U23_MP4$4_source 0 0.0268771f
c_16 U23_MP4$3_source 0 0.0268771f
c_17 U23_MP4$2_source 0 0.0268771f
c_18 U23_MP4$1_source 0 0.0268771f
c_19 U23_MP4$0_source 0 0.0268771f
*
.include "pc3x13.dist.sp.PC3X13.pxi"
*
.ends
*
*
* File: pt3b01d.dist.sp
* Created: Sun Jul  4 12:56:53 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b01d.dist.sp.pex"
.subckt pt3b01d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M56 N_U27_padr_M56_d N_net_m56_VDDO_res_M56_g U28_U22_source N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M57 U28_U22_source N_net_m57_VDDO_res_M57_g N_VSSO_M57_s N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM56 N_net_m56_VDDO_res_RM56_pos N_VDDO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM57 N_VDDO_RM56_neg N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M63 N_U27_padr_M63_d N_net_m63_VSSO_res_M63_g N_VSSO_M63_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M63@2 N_U27_padr_M63@2_d N_net_m63_VSSO_res_M63@2_g N_VSSO_M63_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62 N_U26_MPI1_drain_M62_d N_U27_padr_M62_g N_VSSO_M62_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M64 N_CIN_M64_d N_U26_MPI1_drain_M64_g N_VSS_M64_s N_VSS_M25_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M60 N_U27_padr_M60_d N_net_m60_VDDO_res_M60_g N_VDDO_M60_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 U26_MPI2_drain N_U27_padr_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M59 N_U26_MPI1_drain_M59_d N_U27_padr_M59_g U26_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M61 N_CIN_M61_d N_U26_MPI1_drain_M61_g N_VDD_M61_s N_VDD_M42_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M61@2 N_CIN_M61@2_d N_U26_MPI1_drain_M61@2_g N_VDD_M61_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M61@3 N_CIN_M61@2_d N_U26_MPI1_drain_M61@3_g N_VDD_M61@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M61@4 N_CIN_M61@4_d N_U26_MPI1_drain_M61@4_g N_VDD_M61@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM60 N_net_m60_VDDO_res_RM60_pos N_VDDO_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b01d.dist.sp.PT3B01D.pxi"
*
.ends
*
*
* File: pt3b01.dist.sp
* Created: Sun Jul  4 12:55:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b01.dist.sp.pex"
.subckt pt3b01  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M61 N_U27_padr_M61_d N_net_m61_VSSO_res_M61_g N_VSSO_M61_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M61@2 N_U27_padr_M61@2_d N_net_m61_VSSO_res_M61@2_g N_VSSO_M61_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60 N_U26_MPI1_drain_M60_d N_U27_padr_M60_g N_VSSO_M60_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M62 N_CIN_M62_d N_U26_MPI1_drain_M62_g N_VSS_M62_s N_VSS_M25_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 N_U27_padr_M58_d N_net_m58_VDDO_res_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M56 U26_MPI2_drain N_U27_padr_M56_g N_VDDO_M56_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M57 N_U26_MPI1_drain_M57_d N_U27_padr_M57_g U26_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M59 N_CIN_M59_d N_U26_MPI1_drain_M59_g N_VDD_M59_s N_VDD_M42_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M59@2 N_CIN_M59@2_d N_U26_MPI1_drain_M59@2_g N_VDD_M59_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M59@3 N_CIN_M59@2_d N_U26_MPI1_drain_M59@3_g N_VDD_M59@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M59@4 N_CIN_M59@4_d N_U26_MPI1_drain_M59@4_g N_VDD_M59@3_s N_VDD_M42_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM58 N_net_m58_VDDO_res_RM58_pos N_VDDO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM61 N_VSSO_RM61_pos N_net_m61_VSSO_res_RM61_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b01.dist.sp.PT3B01.pxi"
*
.ends
*
*
* File: pt3b01u.dist.sp
* Created: Sun Jul  4 12:57:03 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b01u.dist.sp.pex"
.subckt pt3b01u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M35 N_PAD_M36_d N_U27_U69$9_gate_M35_g N_VSSO_M35_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U27_U69$9_gate_M36_g N_VSSO_M36_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M37 N_PAD_M38_d N_U27_U69$9_gate_M37_g N_VSSO_M37_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M38_d N_U27_U69$9_gate_M38_g N_VSSO_M35_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M39 N_PAD_M40_d N_U27_U69$9_gate_M39_g N_VSSO_M39_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U27_U69$9_gate_M40_g N_VSSO_M37_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M42_d N_U27_U69$9_gate_M41_g N_VSSO_M41_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M42_d N_U27_U69$9_gate_M42_g N_VSSO_M39_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M43_d N_U15_ngate_M33_g N_VSSO_M33_s N_VSSO_M36_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M43 N_PAD_M43_d N_U27_U69$9_gate_M43_g N_VSSO_M41_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M44 N_PAD_M34_d N_U27_U69$9_gate_M44_g N_VSSO_M44_s N_VSSO_M36_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M34_d N_U15_ngate_M34_g N_VSSO_M33_s N_VSSO_M36_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U27_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M63_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M58 N_U15_pgate_M58_d N_net_m58_VSSO_res_M58_g N_U27_U72_pgate_M58_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M58@2 N_U15_pgate_M58_d N_net_m58_VSSO_res_M58@2_g N_U27_U72_pgate_M58@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@3 N_U15_pgate_M58@3_d N_net_m58_VSSO_res_M58@3_g N_U27_U72_pgate_M58@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@4 N_U15_pgate_M58@3_d N_net_m58_VSSO_res_M58@4_g N_U27_U72_pgate_M58@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M58@5 N_U15_pgate_M58@5_d N_net_m58_VSSO_res_M58@5_g N_U27_U72_pgate_M58@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U27_U69$9_gate_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XR59 N_noxref_2_R59_pos N_PAD_R59_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR60 N_noxref_2_R60_pos N_U27_padr_R60_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M47 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M47_g N_PAD_M47_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M48 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M48_g N_PAD_M47_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M45 N_VDDO_M56_d N_U27_U72_pgate_M45_g N_PAD_M45_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M46 N_VDDO_M46_d N_U27_U72_pgate_M46_g N_PAD_M45_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M49 N_VDDO_M49_d N_U27_U71_UN_P_TOP_M49_g N_PAD_M49_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M50_g N_PAD_M49_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M51 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M51_g N_PAD_M51_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M52_g N_PAD_M51_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M53_g N_PAD_M53_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U27_U71_UN_P_TOP_M54_g N_PAD_M53_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_VDDO_M54_d N_U27_U71_UN_P_TOP_M55_g N_PAD_M55_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M56 N_VDDO_M56_d N_U27_U71_UN_P_TOP_M56_g N_PAD_M55_s N_VDDO_M49_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M57 N_U15_pgate_M57_d N_net_m57_VDDO_res_M57_g N_U27_U72_pgate_M57_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M57@2 N_U15_pgate_M57_d N_net_m57_VDDO_res_M57@2_g N_U27_U72_pgate_M57@2_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M57@3 N_U15_pgate_M57@3_d N_net_m57_VDDO_res_M57@3_g N_U27_U72_pgate_M57@2_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U27_U71_UN_P_TOP_M62_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_U27_padr_M7_d N_net_m7_VSSO_res_M7_g N_VSSO_M7_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M7@2 N_U27_padr_M7@2_d N_net_m7_VSSO_res_M7@2_g N_VSSO_M7_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6 N_U26_MPI1_drain_M6_d N_U27_padr_M6_g N_VSSO_M6_s N_VSS_M57_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M8 N_CIN_M8_d N_U26_MPI1_drain_M8_g N_VSS_M8_s N_VSS_M57_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M30 N_U15_U12_oenb_M30_d N_U15_U15_OUTSHIFT_M30_g N_VSSO_M30_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M9 N_U15_ngate_M9_d N_U15_ISHF_M9_g N_VSSO_M9_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M9@2 N_U15_ngate_M9_d N_U15_ISHF_M9@2_g N_VSSO_M9@2_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M29 N_U15_ngate_M29_d N_U15_U15_OUTSHIFT_M29_g N_VSSO_M9@2_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M10 N_U15_pgate_M10_d N_U15_U12_oenb_M10_g N_U15_ngate_M10_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M10@2 N_U15_pgate_M10@2_d N_U15_U12_oenb_M10@2_g N_U15_ngate_M10_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M10@3 N_U15_pgate_M10@2_d N_U15_U12_oenb_M10@3_g N_U15_ngate_M10@3_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M23 N_U15_U15_MPLL1_dr_M23_d N_OEN_M23_g N_VSSO_M23_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M25 N_VDDO_M25_d N_U15_U15_MN1_drai_M25_g N_U15_U15_MPLL1_dr_M25_s N_VSS_M57_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M23@2 N_U15_U15_MPLL1_dr_M23@2_d N_OEN_M23@2_g N_VSSO_M23_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M24 N_U15_U15_OUTSHIFT_M24_d N_U15_U15_MN1_drai_M24_g N_VSSO_M24_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M24@2 N_U15_U15_OUTSHIFT_M24@2_d N_U15_U15_MN1_drai_M24@2_g N_VSSO_M24_s
+ N_VSS_M57_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M17 N_VDDO_M17_d N_U15_U14_MN1_drai_M17_g N_U15_U14_MPLL1_dr_M17_s N_VSS_M57_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M15 N_U15_U14_MPLL1_dr_M15_d N_I_M15_g N_VSSO_M15_s N_VSS_M57_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M15@2 N_U15_U14_MPLL1_dr_M15@2_d N_I_M15@2_g N_VSSO_M15_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U15_ISHF_M16_d N_U15_U14_MN1_drai_M16_g N_VSSO_M16_s N_VSS_M57_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16@2 N_U15_ISHF_M16@2_d N_U15_U14_MN1_drai_M16@2_g N_VSSO_M16_s N_VSS_M57_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M18 N_U15_U14_MN1_drai_M18_d N_I_M18_g N_VSS_M18_s N_VSS_M57_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M26 N_U15_U15_MN1_drai_M26_d N_OEN_M26_g N_VSS_M18_s N_VSS_M57_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U27_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M4 N_U27_padr_M4_d N_net_m4_VDDO_res_M4_g N_VDDO_M4_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M2 U26_MPI2_drain N_U27_padr_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M3 N_U26_MPI1_drain_M3_d N_U27_padr_M3_g U26_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M31 N_U15_U12_oenb_M31_d N_U15_U15_OUTSHIFT_M31_g N_VDDO_M31_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M31@2 N_U15_U12_oenb_M31@2_d N_U15_U15_OUTSHIFT_M31@2_g N_VDDO_M31_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M11 N_U15_pgate_M11_d N_U15_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M11@2 N_U15_pgate_M11@2_d N_U15_ISHF_M11@2_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M32 N_U15_pgate_M11@2_d N_U15_U12_oenb_M32_g N_VDDO_M32_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M32@2 N_U15_pgate_M32@2_d N_U15_U12_oenb_M32@2_g N_VDDO_M32_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M12 N_U15_ngate_M12_d N_U15_U15_OUTSHIFT_M12_g N_U15_pgate_M12_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M12@2 N_U15_ngate_M12_d N_U15_U15_OUTSHIFT_M12@2_g N_U15_pgate_M12@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M12@3 N_U15_ngate_M12@3_d N_U15_U15_OUTSHIFT_M12@3_g N_U15_pgate_M12@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M21 N_U15_U15_MPLL1_dr_M21_d N_U15_U15_OUTSHIFT_M21_g N_VDDO_M21_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M22 N_U15_U15_OUTSHIFT_M22_d N_U15_U15_MPLL1_dr_M22_g N_VDDO_M21_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M13 N_U15_U14_MPLL1_dr_M13_d N_U15_ISHF_M13_g N_VDDO_M13_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M14 N_U15_ISHF_M14_d N_U15_U14_MPLL1_dr_M14_g N_VDDO_M13_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M5 N_CIN_M5_d N_U26_MPI1_drain_M5_g N_VDD_M5_s N_VDD_M19_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M5@2 N_CIN_M5@2_d N_U26_MPI1_drain_M5@2_g N_VDD_M5_s N_VDD_M19_b PHV L=3.6e-07
+ W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M5@3 N_CIN_M5@2_d N_U26_MPI1_drain_M5@3_g N_VDD_M5@3_s N_VDD_M19_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M5@4 N_CIN_M5@4_d N_U26_MPI1_drain_M5@4_g N_VDD_M5@3_s N_VDD_M19_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M19 N_U15_U14_MN1_drai_M19_d N_I_M19_g N_VDD_M19_s N_VDD_M19_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M19@2 N_U15_U14_MN1_drai_M19_d N_I_M19@2_g N_VDD_M19@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M27 N_U15_U15_MN1_drai_M27_d N_OEN_M27_g N_VDD_M19@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M27@2 N_U15_U15_MN1_drai_M27_d N_OEN_M27@2_g N_VDD_M27@2_s N_VDD_M19_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D20 N_VSS_M57_b N_I_D20_neg DN18  AREA=2.5e-13 PJ=2e-06
D28 N_VSS_M57_b N_OEN_D28_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_net_m4_VDDO_res_RM4_pos N_VDDO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM57 N_VDDO_RM57_pos N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM7 N_VSSO_RM7_pos N_net_m7_VSSO_res_RM7_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM58 N_net_m58_VSSO_res_RM58_pos N_VSSO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b01u.dist.sp.PT3B01U.pxi"
*
.ends
*
*
* File: pt3b02d.dist.sp
* Created: Sun Jul  4 12:58:23 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b02d.dist.sp.pex"
.subckt pt3b02d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M71 N_U28_padr_M71_d N_net_m71_VDDO_res_M71_g U29_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U29_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b02d.dist.sp.PT3B02D.pxi"
*
.ends
*
*
* File: pt3b02.dist.sp
* Created: Sun Jul  4 12:58:19 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b02.dist.sp.pex"
.subckt pt3b02  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b02.dist.sp.PT3B02.pxi"
*
.ends
*
*
* File: pt3b02u.dist.sp
* Created: Sun Jul  4 13:00:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b02u.dist.sp.pex"
.subckt pt3b02u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M71 N_U28_padr_M71_d N_net_m71_VSSO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VSSO_res_RM71_pos N_VSSO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U28_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M31_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U28_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359728f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b02u.dist.sp.PT3B02U.pxi"
*
.ends
*
*
* File: pt3b03d.dist.sp
* Created: Sun Jul  4 13:01:43 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b03d.dist.sp.pex"
.subckt pt3b03d  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M71 N_U29_padr_M71_d N_net_m71_VDDO_res_M71_g U31_U22_source N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M72 U31_U22_source N_net_m72_VDDO_res_M72_g N_VSSO_M72_s N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_net_m71_VDDO_res_RM71_pos N_VDDO_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM72 N_VDDO_RM71_neg N_net_m72_VDDO_res_RM72_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b03d.dist.sp.PT3B03D.pxi"
*
.ends
*
*
* File: pt3b03.dist.sp
* Created: Sun Jul  4 13:00:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b03.dist.sp.pex"
.subckt pt3b03  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b03.dist.sp.PT3B03.pxi"
*
.ends
*
*
* File: pt3b03u.dist.sp
* Created: Sun Jul  4 13:01:49 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3b03u.dist.sp.pex"
.subckt pt3b03u  PAD I OEN CIN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M71 N_U29_padr_M71_d N_net_m71_VSSO_res_M71_g N_VDDO_M71_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM71 N_VSSO_RM71_pos N_net_m71_VSSO_res_RM71_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VSSO_M69_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M69@2 N_U29_padr_M69@2_d N_net_m69_VSSO_res_M69@2_g N_VSSO_M69_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U26_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M70 N_CIN_M70_d N_U26_MPI1_drain_M70_g N_VSS_M70_s N_VSS_M19_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U26_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U26_MPI1_drain_M65_d N_U29_padr_M65_g U26_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M67 N_CIN_M67_d N_U26_MPI1_drain_M67_g N_VDD_M67_s N_VDD_M50_b PHV L=3.6e-07
+ W=8e-06 AD=5.36e-12 AS=3.28e-12 PD=1.734e-05 PS=8.82e-06
M67@2 N_CIN_M67@2_d N_U26_MPI1_drain_M67@2_g N_VDD_M67_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@3 N_CIN_M67@2_d N_U26_MPI1_drain_M67@3_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=3.28e-12 AS=3.28e-12 PD=8.82e-06 PS=8.82e-06
M67@4 N_CIN_M67@4_d N_U26_MPI1_drain_M67@4_g N_VDD_M67@3_s N_VDD_M50_b PHV
+ L=3.6e-07 W=8e-06 AD=4.96e-12 AS=3.28e-12 PD=1.724e-05 PS=8.82e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U26_MPI2_drain 0 0.0169448f
*
.include "pt3b03u.dist.sp.PT3B03U.pxi"
*
.ends
*
*
* File: pt3o01.dist.sp
* Created: Sun Jul  4 13:03:17 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3o01.dist.sp.pex"
.subckt pt3o01  PAD I VDD VSS VDDO VSSO 
* 
M29 N_ngate_M29_d N_U28_ISHF_M29_g N_VSSO_M29_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M29@2 N_ngate_M29_d N_U28_ISHF_M29@2_g N_VSSO_M29@2_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.6e-12 PD=1.082e-05 PS=2.132e-05
M30 N_pgate_M30_d N_net_m30_VDDO_res_M30_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M30@2 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@2_g N_ngate_M30_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M30@3 N_pgate_M30@2_d N_net_m30_VDDO_res_M30@3_g N_ngate_M30@3_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M37 N_VDDO_M37_d N_U28_U16_MN1_drai_M37_g N_U28_U16_MPLL1_dr_M37_s N_VSS_M29_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M35 N_U28_U16_MPLL1_dr_M35_d N_I_M35_g N_VSSO_M35_s N_VSS_M29_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M35@2 N_U28_U16_MPLL1_dr_M35@2_d N_I_M35@2_g N_VSSO_M35_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36 N_U28_ISHF_M36_d N_U28_U16_MN1_drai_M36_g N_VSSO_M36_s N_VSS_M29_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M36@2 N_U28_ISHF_M36@2_d N_U28_U16_MN1_drai_M36@2_g N_VSSO_M36_s N_VSS_M29_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5 N_PAD_M11_d N_U29_U74$9_gate_M5_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M12_d N_U29_U74$9_gate_M6_g N_VSSO_M6_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M13_d N_U29_U74$9_gate_M7_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M14_d N_U29_U74$9_gate_M8_g N_VSSO_M5_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M3_d N_U29_U74$9_gate_M9_g N_VSSO_M9_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M4_d N_U29_U74$9_gate_M10_g N_VSSO_M7_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_U28_U16_MN1_drai_M38_d N_I_M38_g N_VSS_M38_s N_VSS_M29_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M31 N_pgate_M31_d N_U28_ISHF_M31_g N_VDDO_M31_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.32e-11 AS=8.2e-12 PD=4.132e-05 PS=2.082e-05
M31@2 N_pgate_M31@2_d N_U28_ISHF_M31@2_g N_VDDO_M31_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M32 N_ngate_M32_d N_net_m32_VSSO_res_M32_g N_pgate_M32_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_ngate_M32_d N_net_m32_VSSO_res_M32@2_g N_pgate_M32@2_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M32@3 N_ngate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_pgate_M32@2_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33 N_U28_U16_MPLL1_dr_M33_d N_U28_ISHF_M33_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M34 N_U28_ISHF_M34_d N_U28_U16_MPLL1_dr_M34_g N_VDDO_M33_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M39 N_U28_U16_MN1_drai_M39_d N_I_M39_g N_VDD_M39_s N_VDD_M39_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M39@2 N_U28_U16_MN1_drai_M39_d N_I_M39@2_g N_VDD_M39@2_s N_VDD_M39_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D40 N_VSS_M29_b N_I_D40_neg DN18  AREA=2.5e-13 PJ=2e-06
XR27 N_VSSO_R27_pos N_U29_U74$9_gate_R27_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR28 N_U29_U37_r2_R28_pos N_VDDO_R28_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M11 N_PAD_M11_d N_U29_U74$9_gate_M11_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_U74$9_gate_M12_g N_VSSO_M11_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U74$9_gate_M13_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U29_U74$9_gate_M14_g N_VSSO_M13_s N_VSSO_M11_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M3 N_PAD_M3_d N_ngate_M3_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_ngate_M4_g N_VSSO_M3_s N_VSSO_M11_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR1 U29_U69_padr N_noxref_11_R1_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR2 N_noxref_11_R2_pos N_PAD_R2_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XRM30 N_net_m30_VDDO_res_RM30_pos N_VDDO_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
M17 N_VDDO_M17_d N_U29_U37_r2_M17_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M18 N_VDDO_M19_d N_U29_U37_r2_M18_g N_PAD_M17_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M15 N_VDDO_M26_d N_pgate_M15_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M16 N_VDDO_M16_d N_pgate_M16_g N_PAD_M15_s N_VDDO_M19_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M19 N_VDDO_M19_d N_U29_U37_r2_M19_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U29_U37_r2_M20_g N_PAD_M19_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U29_U37_r2_M21_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U29_U37_r2_M22_g N_PAD_M21_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U29_U37_r2_M23_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U29_U37_r2_M24_g N_PAD_M23_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M24_d N_U29_U37_r2_M25_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U37_r2_M26_g N_PAD_M25_s N_VDDO_M19_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
c_1 U29_U69_padr 0 17.4974f
*
.include "pt3o01.dist.sp.PT3O01.pxi"
*
.ends
*
*
* File: pt3o02.dist.sp
* Created: Sun Jul  4 13:03:24 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3o02.dist.sp.pex"
.subckt pt3o02  PAD I VDD VSS VDDO VSSO 
* 
M13 N_PAD_M17_d N_U29_U76_r1_M13_g N_VSSO_M13_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M18_d N_U29_U76_r1_M14_g N_VSSO_M14_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M9 N_PAD_M7_d N_U30_ngate2_M9_g N_VSSO_M9_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M15 N_PAD_M8_d N_U29_U76_r1_M15_g N_VSSO_M13_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M11_d N_U29_U76_r1_M16_g N_VSSO_M16_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M12_d N_U30_ngate2_M10_g N_VSSO_M9_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M17 N_PAD_M17_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U29_U76_r1_M18_g N_VSSO_M17_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M7_d N_ngate_M7_g N_VSSO_M7_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_ngate_M8_g N_VSSO_M7_s N_VSSO_M17_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U29_ngate3_M11_g N_VSSO_M11_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_ngate3_M12_g N_VSSO_M11_s N_VSSO_M17_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR31 U29_U69_padr N_noxref_2_R31_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR32 N_noxref_2_R32_pos N_PAD_R32_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U29_U37_r2_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U29_U37_r2_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U37_r2_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U37_r2_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U37_r2_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U37_r2_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M34 N_U29_ngate3_M34_d N_U30_ngatex_M34_g N_VSSO_M34_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U28_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U28_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U28_U13_MN1_drai_M45_g N_U28_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U28_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U28_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U28_ISHF_M44_d N_U28_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U28_ISHF_M44@2_d N_U28_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U28_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M33 N_U29_ngate3_M33_d N_U30_ngatex_M33_g N_U30_ngate2_M33_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U28_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U28_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U28_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U28_U13_MPLL1_dr_M41_d N_U28_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U28_ISHF_M42_d N_U28_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U28_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U28_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.5122f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pt3o02.dist.sp.PT3O02.pxi"
*
.ends
*
*
* File: pt3o03.dist.sp
* Created: Sun Jul  4 13:05:17 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3o03.dist.sp.pex"
.subckt pt3o03  PAD I VDD VSS VDDO VSSO 
* 
M13 N_PAD_M15_d N_ngate_M13_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M16_d N_U29_U76_r1_M17_g N_VSSO_M17_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M7 N_PAD_M9_d N_U30_ngate2_M7_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M10_d N_ngate_M14_g N_VSSO_M13_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M11_d N_U29_U76_r1_M18_g N_VSSO_M18_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M12_d N_U30_ngate2_M8_g N_VSSO_M7_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR35 N_VSSO_R35_pos N_U29_U76_r1_R35_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR36 N_U29_U37_r2_R36_pos N_VDDO_R36_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
M15 N_PAD_M15_d N_ngate_M15_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_ngate_M16_g N_VSSO_M15_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M9_d N_U30_ngate2_M9_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U30_ngate2_M10_g N_VSSO_M9_s N_VSSO_M15_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U29_ngate3_M11_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U29_ngate3_M12_g N_VSSO_M11_s N_VSSO_M15_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
XR19 U29_U69_padr N_noxref_2_R19_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR20 N_noxref_2_R20_pos N_PAD_R20_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M33 N_VDDO_M33_d N_U29_U37_r2_M33_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M34 N_VDDO_M25_d N_U29_U37_r2_M34_g N_PAD_M33_s N_VDDO_M25_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M32_d N_pgate_M23_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_pgate_M24_g N_PAD_M23_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M25 N_VDDO_M25_d N_pgate_M25_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_pgate_M26_g N_PAD_M25_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M27 N_VDDO_M26_d N_pgate_M27_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_pgate_M28_g N_PAD_M27_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_pgate_M29_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_pgate_M30_g N_PAD_M29_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_pgate_M31_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_pgate_M32_g N_PAD_M31_s N_VDDO_M25_b PHV L=4e-07 W=5.2e-05
+ AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M3 N_U30_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M3_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U30_ngate2_M4_d N_U30_ngatex_M4_g N_VSSO_M4_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U30_ngatex_M1_d N_ngate_M1_g N_VSSO_M1_s N_VSS_M3_b NHV L=3.6e-07 W=1e-05
+ AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M22 N_U29_ngate3_M22_d N_U30_ngatex_M22_g N_VSSO_M22_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M39 N_ngate_M39_d N_U27_ISHF_M39_g N_VSSO_M39_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M39@2 N_ngate_M39_d N_U27_ISHF_M39@2_g N_VSSO_M39@2_s N_VSS_M3_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M40 N_pgate_M40_d N_net_m40_VDDO_res_M40_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M40@2 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@2_g N_ngate_M40_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M40@3 N_pgate_M40@2_d N_net_m40_VDDO_res_M40@3_g N_ngate_M40@3_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M45 N_VDDO_M45_d N_U27_U13_MN1_drai_M45_g N_U27_U13_MPLL1_dr_M45_s N_VSS_M3_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M43 N_U27_U13_MPLL1_dr_M43_d N_I_M43_g N_VSSO_M43_s N_VSS_M3_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U27_U13_MPLL1_dr_M43@2_d N_I_M43@2_g N_VSSO_M43_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44 N_U27_ISHF_M44_d N_U27_U13_MN1_drai_M44_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M44@2 N_U27_ISHF_M44@2_d N_U27_U13_MN1_drai_M44@2_g N_VSSO_M44_s N_VSS_M3_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46 N_U27_U13_MN1_drai_M46_d N_I_M46_g N_VSS_M46_s N_VSS_M3_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=2.925e-12 PD=1.117e-05 PS=1.117e-05
M6 U30_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M6_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U30_ngate2_M5_d N_U30_ngatex_M5_g U30_U15_U8_sourc N_VDDO_M6_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U30_ngatex_M2_d N_ngate_M2_g N_VDDO_M2_s N_VDDO_M6_b PHV L=3.6e-07 W=7e-06
+ AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M21 N_U29_ngate3_M21_d N_U30_ngatex_M21_g N_U30_ngate2_M21_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M37 N_pgate_M37_d N_U27_ISHF_M37_g N_VDDO_M37_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M37@2 N_pgate_M37_d N_U27_ISHF_M37@2_g N_VDDO_M37@2_s N_VDDO_M6_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M37@3 N_pgate_M37@3_d N_U27_ISHF_M37@3_g N_VDDO_M37@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=8.2e-12 PD=4.124e-05 PS=2.082e-05
M38 N_ngate_M38_d N_net_m38_VSSO_res_M38_g N_pgate_M38_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M38@2 N_ngate_M38_d N_net_m38_VSSO_res_M38@2_g N_pgate_M38@2_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M38@3 N_ngate_M38@3_d N_net_m38_VSSO_res_M38@3_g N_pgate_M38@2_s N_VDDO_M6_b
+ PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05 PS=1.082e-05
M41 N_U27_U13_MPLL1_dr_M41_d N_U27_ISHF_M41_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U27_ISHF_M42_d N_U27_U13_MPLL1_dr_M42_g N_VDDO_M41_s N_VDDO_M6_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M47 N_U27_U13_MN1_drai_M47_d N_I_M47_g N_VDD_M47_s N_VDD_M47_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M47@2 N_U27_U13_MN1_drai_M47_d N_I_M47@2_g N_VDD_M47@2_s N_VDD_M47_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=3.1e-12 PD=5.56e-06 PS=1.124e-05
D48 N_VSS_M3_b N_I_D48_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM40 N_net_m40_VDDO_res_RM40_pos N_VDDO_RM40_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_net_m38_VSSO_res_RM38_pos N_VSSO_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_U69_padr 0 17.4884f
c_2 U30_U15_U8_sourc 0 0.360661f
*
.include "pt3o03.dist.sp.PT3O03.pxi"
*
.ends
*
*
* File: pt3t01d.dist.sp
* Created: Sun Jul  4 13:06:52 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t01d.dist.sp.pex"
.subckt pt3t01d  PAD I OEN VDD VSS VDDO VSSO 
* 
M56 N_U27_padr_M56_d N_net_m56_VDDO_res_M56_g U28_U22_source N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M57 U28_U22_source N_net_m57_VDDO_res_M57_g N_VSSO_M57_s N_VSS_M25_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM56 N_net_m56_VDDO_res_RM56_pos N_VDDO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM57 N_VDDO_RM56_neg N_net_m57_VDDO_res_RM57_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M61 N_U27_padr_M61_d N_net_m61_VSSO_res_M61_g N_VSSO_M61_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M61@2 N_U27_padr_M61@2_d N_net_m61_VSSO_res_M61@2_g N_VSSO_M61_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62 N_U29_MPI1_drain_M62_d N_U27_padr_M62_g N_VSSO_M62_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M60 N_U27_padr_M60_d N_net_m60_VDDO_res_M60_g N_VDDO_M60_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 U29_MPI2_drain N_U27_padr_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M59 N_U29_MPI1_drain_M59_d N_U27_padr_M59_g U29_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM60 N_net_m60_VDDO_res_RM60_pos N_VDDO_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM61 N_VSSO_RM61_pos N_net_m61_VSSO_res_RM61_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_MPI2_drain 0 0.0289375f
*
.include "pt3t01d.dist.sp.PT3T01D.pxi"
*
.ends
*
*
* File: pt3t01.dist.sp
* Created: Sun Jul  4 13:05:03 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t01.dist.sp.pex"
.subckt pt3t01  PAD I OEN VDD VSS VDDO VSSO 
* 
M3 N_PAD_M4_d N_U27_U69$9_gate_M3_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M4 N_PAD_M4_d N_U27_U69$9_gate_M4_g N_VSSO_M4_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M5 N_PAD_M6_d N_U27_U69$9_gate_M5_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M6 N_PAD_M6_d N_U27_U69$9_gate_M6_g N_VSSO_M3_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M8_d N_U27_U69$9_gate_M7_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U27_U69$9_gate_M8_g N_VSSO_M5_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M10_d N_U27_U69$9_gate_M9_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M10_d N_U27_U69$9_gate_M10_g N_VSSO_M7_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_PAD_M11_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U27_U69$9_gate_M11_g N_VSSO_M9_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M2_d N_U27_U69$9_gate_M12_g N_VSSO_M12_s N_VSSO_M4_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M2 N_PAD_M2_d N_U15_ngate_M2_g N_VSSO_M1_s N_VSSO_M4_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M26 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26_g N_U27_U72_pgate_M26_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M26@2 N_U15_pgate_M26_d N_net_m26_VSSO_res_M26@2_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@3 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@3_g N_U27_U72_pgate_M26@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@4 N_U15_pgate_M26@3_d N_net_m26_VSSO_res_M26@4_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M26@5 N_U15_pgate_M26@5_d N_net_m26_VSSO_res_M26@5_g N_U27_U72_pgate_M26@4_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR29 N_U27_U69$9_gate_R29_pos N_VSSO_R29_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR27 N_noxref_2_R27_pos N_PAD_R27_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR28 N_noxref_2_R28_pos N_U27_padr_R28_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M15 N_VDDO_M15_d N_U27_U71_UN_P_TOP_M15_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M16 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M16_g N_PAD_M15_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M13 N_VDDO_M24_d N_U27_U72_pgate_M13_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M14 N_VDDO_M14_d N_U27_U72_pgate_M14_g N_PAD_M13_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M17 N_VDDO_M17_d N_U27_U71_UN_P_TOP_M17_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M18 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M18_g N_PAD_M17_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M18_d N_U27_U71_UN_P_TOP_M19_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M20_g N_PAD_M19_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M20_d N_U27_U71_UN_P_TOP_M21_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M22_g N_PAD_M21_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U27_U71_UN_P_TOP_M23_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U27_U71_UN_P_TOP_M24_g N_PAD_M23_s N_VDDO_M17_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25_g N_U27_U72_pgate_M25_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M25@2 N_U15_pgate_M25_d N_net_m25_VDDO_res_M25@2_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M25@3 N_U15_pgate_M25@3_d N_net_m25_VDDO_res_M25@3_g N_U27_U72_pgate_M25@2_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M30 N_VDDO_M30_d N_net_m30_VDDO_res_M30_g N_U27_U71_UN_P_TOP_M30_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M59 N_U27_padr_M59_d N_net_m59_VSSO_res_M59_g N_VSSO_M59_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M59@2 N_U27_padr_M59@2_d N_net_m59_VSSO_res_M59@2_g N_VSSO_M59_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M60 N_U28_MPI1_drain_M60_d N_U27_padr_M60_g N_VSSO_M60_s N_VSS_M25_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M53 N_U15_U12_oenb_M53_d N_U15_U15_OUTSHIFT_M53_g N_VSSO_M53_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M32 N_U15_ngate_M32_d N_U15_ISHF_M32_g N_VSSO_M32_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M32@2 N_U15_ngate_M32_d N_U15_ISHF_M32@2_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M52 N_U15_ngate_M52_d N_U15_U15_OUTSHIFT_M52_g N_VSSO_M32@2_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M33 N_U15_pgate_M33_d N_U15_U12_oenb_M33_g N_U15_ngate_M33_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M33@2 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@2_g N_U15_ngate_M33_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M33@3 N_U15_pgate_M33@2_d N_U15_U12_oenb_M33@3_g N_U15_ngate_M33@3_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M46 N_U15_U15_MPLL1_dr_M46_d N_OEN_M46_g N_VSSO_M46_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U15_MN1_drai_M48_g N_U15_U15_MPLL1_dr_M48_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46@2 N_U15_U15_MPLL1_dr_M46@2_d N_OEN_M46@2_g N_VSSO_M46_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_U15_OUTSHIFT_M47_d N_U15_U15_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_U15_OUTSHIFT_M47@2_d N_U15_U15_MN1_drai_M47@2_g N_VSSO_M47_s
+ N_VSS_M25_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_VDDO_M40_d N_U15_U14_MN1_drai_M40_g N_U15_U14_MPLL1_dr_M40_s N_VSS_M25_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M38 N_U15_U14_MPLL1_dr_M38_d N_I_M38_g N_VSSO_M38_s N_VSS_M25_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M38@2 N_U15_U14_MPLL1_dr_M38@2_d N_I_M38@2_g N_VSSO_M38_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39 N_U15_ISHF_M39_d N_U15_U14_MN1_drai_M39_g N_VSSO_M39_s N_VSS_M25_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M39@2 N_U15_ISHF_M39@2_d N_U15_U14_MN1_drai_M39@2_g N_VSSO_M39_s N_VSS_M25_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U15_U14_MN1_drai_M41_d N_I_M41_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M49 N_U15_U15_MN1_drai_M49_d N_OEN_M49_g N_VSS_M41_s N_VSS_M25_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M31 N_U27_U71_UN_P_TOP_M31_d N_net_m31_VSSO_res_M31_g N_VDDO_M31_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M58 N_U27_padr_M58_d N_net_m58_VDDO_res_M58_g N_VDDO_M58_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M56 U28_MPI2_drain N_U27_padr_M56_g N_VDDO_M56_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M57 N_U28_MPI1_drain_M57_d N_U27_padr_M57_g U28_MPI2_drain N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M54 N_U15_U12_oenb_M54_d N_U15_U15_OUTSHIFT_M54_g N_VDDO_M54_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M54@2 N_U15_U12_oenb_M54@2_d N_U15_U15_OUTSHIFT_M54@2_g N_VDDO_M54_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M34 N_U15_pgate_M34_d N_U15_ISHF_M34_g N_VDDO_M34_s N_VDDO_M31_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M34@2 N_U15_pgate_M34@2_d N_U15_ISHF_M34@2_g N_VDDO_M34_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M55 N_U15_pgate_M34@2_d N_U15_U12_oenb_M55_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M55@2 N_U15_pgate_M55@2_d N_U15_U12_oenb_M55@2_g N_VDDO_M55_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M35 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35_g N_U15_pgate_M35_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M35@2 N_U15_ngate_M35_d N_U15_U15_OUTSHIFT_M35@2_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M35@3 N_U15_ngate_M35@3_d N_U15_U15_OUTSHIFT_M35@3_g N_U15_pgate_M35@2_s
+ N_VDDO_M31_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M44 N_U15_U15_MPLL1_dr_M44_d N_U15_U15_OUTSHIFT_M44_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_U15_OUTSHIFT_M45_d N_U15_U15_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M31_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M36 N_U15_U14_MPLL1_dr_M36_d N_U15_ISHF_M36_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M37 N_U15_ISHF_M37_d N_U15_U14_MPLL1_dr_M37_g N_VDDO_M36_s N_VDDO_M31_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M42 N_U15_U14_MN1_drai_M42_d N_I_M42_g N_VDD_M42_s N_VDD_M42_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M42@2 N_U15_U14_MN1_drai_M42_d N_I_M42@2_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50 N_U15_U15_MN1_drai_M50_d N_OEN_M50_g N_VDD_M42@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M50@2 N_U15_U15_MN1_drai_M50_d N_OEN_M50@2_g N_VDD_M50@2_s N_VDD_M42_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D43 N_VSS_M25_b N_I_D43_neg DN18  AREA=2.5e-13 PJ=2e-06
D51 N_VSS_M25_b N_OEN_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM31 N_VSSO_RM31_pos N_net_m31_VSSO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM58 N_net_m58_VDDO_res_RM58_pos N_VDDO_RM58_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM25 N_VDDO_RM25_pos N_net_m25_VDDO_res_RM25_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM30 N_VDDO_RM30_pos N_net_m30_VDDO_res_RM30_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM59 N_VSSO_RM59_pos N_net_m59_VSSO_res_RM59_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM26 N_net_m26_VSSO_res_RM26_pos N_VSSO_RM26_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U28_MPI2_drain 0 0.0289375f
*
.include "pt3t01.dist.sp.PT3T01.pxi"
*
.ends
*
*
* File: pt3t01u.dist.sp
* Created: Sun Jul  4 13:06:37 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t01u.dist.sp.pex"
.subckt pt3t01u  PAD I OEN VDD VSS VDDO VSSO 
* 
M33 N_PAD_M34_d N_U27_U69$9_gate_M33_g N_VSSO_M33_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M34 N_PAD_M34_d N_U27_U69$9_gate_M34_g N_VSSO_M34_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M35 N_PAD_M36_d N_U27_U69$9_gate_M35_g N_VSSO_M35_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U27_U69$9_gate_M36_g N_VSSO_M33_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M37 N_PAD_M38_d N_U27_U69$9_gate_M37_g N_VSSO_M37_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M38_d N_U27_U69$9_gate_M38_g N_VSSO_M35_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M39 N_PAD_M40_d N_U27_U69$9_gate_M39_g N_VSSO_M39_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U27_U69$9_gate_M40_g N_VSSO_M37_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M31 N_PAD_M41_d N_U15_ngate_M31_g N_VSSO_M31_s N_VSSO_M34_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M41_d N_U27_U69$9_gate_M41_g N_VSSO_M39_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M32_d N_U27_U69$9_gate_M42_g N_VSSO_M42_s N_VSSO_M34_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M32 N_PAD_M32_d N_U15_ngate_M32_g N_VSSO_M31_s N_VSSO_M34_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M1 N_U27_padr_M1_d N_net_m1_VSSO_res_M1_g N_VDDO_M1_s N_VDDO_M61_b PHV L=2e-06
+ W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M56 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56_g N_U27_U72_pgate_M56_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M56@2 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56@2_g N_U27_U72_pgate_M56@2_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@3 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@3_g N_U27_U72_pgate_M56@2_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@4 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@4_g N_U27_U72_pgate_M56@4_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@5 N_U15_pgate_M56@5_d N_net_m56_VSSO_res_M56@5_g N_U27_U72_pgate_M56@4_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR59 N_U27_U69$9_gate_R59_pos N_VSSO_R59_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM1 N_net_m1_VSSO_res_RM1_pos N_VSSO_RM1_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XR57 N_noxref_2_R57_pos N_PAD_R57_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR58 N_noxref_2_R58_pos N_U27_padr_R58_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M45 N_VDDO_M45_d N_U27_U71_UN_P_TOP_M45_g N_PAD_M45_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M46 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M46_g N_PAD_M45_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M54_d N_U27_U72_pgate_M43_g N_PAD_M43_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M44 N_VDDO_M44_d N_U27_U72_pgate_M44_g N_PAD_M43_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M47 N_VDDO_M47_d N_U27_U71_UN_P_TOP_M47_g N_PAD_M47_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M48 N_VDDO_M48_d N_U27_U71_UN_P_TOP_M48_g N_PAD_M47_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M49 N_VDDO_M48_d N_U27_U71_UN_P_TOP_M49_g N_PAD_M49_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M50 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M50_g N_PAD_M49_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M51 N_VDDO_M50_d N_U27_U71_UN_P_TOP_M51_g N_PAD_M51_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M52_g N_PAD_M51_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U27_U71_UN_P_TOP_M53_g N_PAD_M53_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U27_U71_UN_P_TOP_M54_g N_PAD_M53_s N_VDDO_M47_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55_g N_U27_U72_pgate_M55_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M55@2 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55@2_g N_U27_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M55@3 N_U15_pgate_M55@3_d N_net_m55_VDDO_res_M55@3_g N_U27_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M60 N_VDDO_M60_d N_net_m60_VDDO_res_M60_g N_U27_U71_UN_P_TOP_M60_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M5 N_U27_padr_M5_d N_net_m5_VSSO_res_M5_g N_VSSO_M5_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M5@2 N_U27_padr_M5@2_d N_net_m5_VSSO_res_M5@2_g N_VSSO_M5_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M6 N_U29_MPI1_drain_M6_d N_U27_padr_M6_g N_VSSO_M6_s N_VSS_M55_b NHV L=3.6e-07
+ W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M28 N_U15_U12_oenb_M28_d N_U15_U15_OUTSHIFT_M28_g N_VSSO_M28_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_U15_ngate_M7_d N_U15_ISHF_M7_g N_VSSO_M7_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M7@2 N_U15_ngate_M7_d N_U15_ISHF_M7@2_g N_VSSO_M7@2_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M27 N_U15_ngate_M27_d N_U15_U15_OUTSHIFT_M27_g N_VSSO_M7@2_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M8 N_U15_pgate_M8_d N_U15_U12_oenb_M8_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@2_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@3_g N_U15_ngate_M8@3_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M21 N_U15_U15_MPLL1_dr_M21_d N_OEN_M21_g N_VSSO_M21_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M23 N_VDDO_M23_d N_U15_U15_MN1_drai_M23_g N_U15_U15_MPLL1_dr_M23_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M21@2 N_U15_U15_MPLL1_dr_M21@2_d N_OEN_M21@2_g N_VSSO_M21_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22 N_U15_U15_OUTSHIFT_M22_d N_U15_U15_MN1_drai_M22_g N_VSSO_M22_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22@2 N_U15_U15_OUTSHIFT_M22@2_d N_U15_U15_MN1_drai_M22@2_g N_VSSO_M22_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M15 N_VDDO_M15_d N_U15_U14_MN1_drai_M15_g N_U15_U14_MPLL1_dr_M15_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U15_U14_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U15_U14_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U15_ISHF_M14_d N_U15_U14_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U15_ISHF_M14@2_d N_U15_U14_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U15_U14_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M24 N_U15_U15_MN1_drai_M24_d N_OEN_M24_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M61 N_U27_U71_UN_P_TOP_M61_d N_net_m61_VSSO_res_M61_g N_VDDO_M61_s N_VDDO_M61_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M4 N_U27_padr_M4_d N_net_m4_VDDO_res_M4_g N_VDDO_M4_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M2 U29_MPI2_drain N_U27_padr_M2_g N_VDDO_M2_s N_VDDO_M61_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M3 N_U29_MPI1_drain_M3_d N_U27_padr_M3_g U29_MPI2_drain N_VDDO_M61_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M29 N_U15_U12_oenb_M29_d N_U15_U15_OUTSHIFT_M29_g N_VDDO_M29_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M29@2 N_U15_U12_oenb_M29@2_d N_U15_U15_OUTSHIFT_M29@2_g N_VDDO_M29_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M9 N_U15_pgate_M9_d N_U15_ISHF_M9_g N_VDDO_M9_s N_VDDO_M61_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M9@2 N_U15_pgate_M9@2_d N_U15_ISHF_M9@2_g N_VDDO_M9_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M30 N_U15_pgate_M9@2_d N_U15_U12_oenb_M30_g N_VDDO_M30_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M30@2 N_U15_pgate_M30@2_d N_U15_U12_oenb_M30@2_g N_VDDO_M30_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M10 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10_g N_U15_pgate_M10_s N_VDDO_M61_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M10@2 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10@2_g N_U15_pgate_M10@2_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M10@3 N_U15_ngate_M10@3_d N_U15_U15_OUTSHIFT_M10@3_g N_U15_pgate_M10@2_s
+ N_VDDO_M61_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M19 N_U15_U15_MPLL1_dr_M19_d N_U15_U15_OUTSHIFT_M19_g N_VDDO_M19_s N_VDDO_M61_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M20 N_U15_U15_OUTSHIFT_M20_d N_U15_U15_MPLL1_dr_M20_g N_VDDO_M19_s N_VDDO_M61_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U15_U14_MPLL1_dr_M11_d N_U15_ISHF_M11_g N_VDDO_M11_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U15_ISHF_M12_d N_U15_U14_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M61_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M17 N_U15_U14_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U15_U14_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25 N_U15_U15_MN1_drai_M25_d N_OEN_M25_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25@2 N_U15_U15_MN1_drai_M25_d N_OEN_M25@2_g N_VDD_M25@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D18 N_VSS_M55_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
D26 N_VSS_M55_b N_OEN_D26_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM61 N_VSSO_RM61_pos N_net_m61_VSSO_res_RM61_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM4 N_net_m4_VDDO_res_RM4_pos N_VDDO_RM4_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM55 N_VDDO_RM55_pos N_net_m55_VDDO_res_RM55_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM60 N_VDDO_RM60_pos N_net_m60_VDDO_res_RM60_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM5 N_VSSO_RM5_pos N_net_m5_VSSO_res_RM5_neg RPMPOLY2T w=2e-06 l=6.455e-06 
XRM56 N_net_m56_VSSO_res_RM56_pos N_VSSO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U29_MPI2_drain 0 0.0289375f
*
.include "pt3t01u.dist.sp.PT3T01U.pxi"
*
.ends
*
*
* File: pt3t02d.dist.sp
* Created: Sun Jul  4 13:08:16 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t02d.dist.sp.pex"
.subckt pt3t02d  PAD I OEN VDD VSS VDDO VSSO 
* 
M69 N_U28_padr_M69_d N_net_m69_VDDO_res_M69_g U29_U22_source N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U29_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M31_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pt3t02d.dist.sp.PT3T02D.pxi"
*
.ends
*
*
* File: pt3t02.dist.sp
* Created: Sun Jul  4 13:08:13 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t02.dist.sp.pex"
.subckt pt3t02  PAD I OEN VDD VSS VDDO VSSO 
* 
M13 N_PAD_M14_d N_U28_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M14_d N_U28_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M15 N_PAD_M16_d N_U28_U42_r1_M15_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M16 N_PAD_M16_d N_U28_U42_r1_M16_g N_VSSO_M13_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M17_d N_U15_ngate_M11_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U28_U42_r1_M17_g N_VSSO_M15_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U17_ngate2_M7_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U15_ngate_M12_g N_VSSO_M11_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M8_d N_U28_ngate3_M9_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M8 N_PAD_M8_d N_U17_ngate2_M8_g N_VSSO_M7_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M10_d N_U28_U42_r1_M18_g N_VSSO_M18_s N_VSSO_M14_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M10 N_PAD_M10_d N_U28_ngate3_M10_g N_VSSO_M9_s N_VSSO_M14_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32_g N_U28_U72_pgate_M32_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M32@2 N_U15_pgate_M32_d N_net_m32_VSSO_res_M32@2_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@3 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@3_g N_U28_U72_pgate_M32@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@4 N_U15_pgate_M32@3_d N_net_m32_VSSO_res_M32@4_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M32@5 N_U15_pgate_M32@5_d N_net_m32_VSSO_res_M32@5_g N_U28_U72_pgate_M32@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U28_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR33 N_noxref_2_R33_pos N_PAD_R33_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR34 N_noxref_2_R34_pos N_U28_padr_R34_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M25 N_VDDO_M25_d N_U28_U71_UN_P_TOP_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M26 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_VDDO_M24_d N_U28_U72_pgate_M19_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M20 N_VDDO_M20_d N_U28_U72_pgate_M20_g N_PAD_M19_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U28_U71_UN_P_TOP_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U28_U71_UN_P_TOP_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U28_U71_UN_P_TOP_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M21 N_VDDO_M30_d N_U28_U72_pgate_M21_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M22 N_VDDO_M22_d N_U28_U72_pgate_M22_g N_PAD_M21_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M23 N_VDDO_M22_d N_U28_U72_pgate_M23_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M24 N_VDDO_M24_d N_U28_U72_pgate_M24_g N_PAD_M23_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31_g N_U28_U72_pgate_M31_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M31@2 N_U15_pgate_M31_d N_net_m31_VDDO_res_M31@2_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M31@3 N_U15_pgate_M31@3_d N_net_m31_VDDO_res_M31@3_g N_U28_U72_pgate_M31@2_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U28_U71_UN_P_TOP_M38_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M31_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M36 N_U28_ngate3_M36_d N_U17_ngatex_M36_g N_VSSO_M36_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M31_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U15_U12_oenb_M61_d N_U15_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M40 N_U15_ngate_M40_d N_U15_ISHF_M40_g N_VSSO_M40_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M40@2 N_U15_ngate_M40_d N_U15_ISHF_M40@2_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M60 N_U15_ngate_M60_d N_U15_U15_OUTSHIFT_M60_g N_VSSO_M40@2_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M41 N_U15_pgate_M41_d N_U15_U12_oenb_M41_g N_U15_ngate_M41_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41@2 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@2_g N_U15_ngate_M41_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M41@3 N_U15_pgate_M41@2_d N_U15_U12_oenb_M41@3_g N_U15_ngate_M41@3_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U15_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U15_U15_MN1_drai_M56_g N_U15_U15_MPLL1_dr_M56_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U15_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U15_U15_OUTSHIFT_M55_d N_U15_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U15_U15_OUTSHIFT_M55@2_d N_U15_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M31_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U15_U14_MN1_drai_M48_g N_U15_U14_MPLL1_dr_M48_s N_VSS_M31_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U15_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M31_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U15_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U15_ISHF_M47_d N_U15_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M31_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U15_ISHF_M47@2_d N_U15_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M31_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U15_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U15_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M31_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U28_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M35 N_U28_ngate3_M35_d N_U17_ngatex_M35_g N_U17_ngate2_M35_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U15_U12_oenb_M62_d N_U15_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U15_U12_oenb_M62@2_d N_U15_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M42 N_U15_pgate_M42_d N_U15_ISHF_M42_g N_VDDO_M42_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M42@2 N_U15_pgate_M42@2_d N_U15_ISHF_M42@2_g N_VDDO_M42_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U15_pgate_M42@2_d N_U15_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U15_pgate_M63@2_d N_U15_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M43 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43_g N_U15_pgate_M43_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M43@2 N_U15_ngate_M43_d N_U15_U15_OUTSHIFT_M43@2_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M43@3 N_U15_ngate_M43@3_d N_U15_U15_OUTSHIFT_M43@3_g N_U15_pgate_M43@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M52 N_U15_U15_MPLL1_dr_M52_d N_U15_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U15_U15_OUTSHIFT_M53_d N_U15_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U15_U14_MPLL1_dr_M44_d N_U15_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U15_ISHF_M45_d N_U15_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U15_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U15_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U15_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U15_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M31_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M31_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM31 N_VDDO_RM31_pos N_net_m31_VDDO_res_RM31_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM32 N_net_m32_VSSO_res_RM32_pos N_VSSO_RM32_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pt3t02.dist.sp.PT3T02.pxi"
*
.ends
*
*
* File: pt3t02u.dist.sp
* Created: Sun Jul  4 13:09:56 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t02u.dist.sp.pex"
.subckt pt3t02u  PAD I OEN VDD VSS VDDO VSSO 
* 
M37 N_PAD_M38_d N_U28_U42_r1_M37_g N_VSSO_M37_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M38 N_PAD_M38_d N_U28_U42_r1_M38_g N_VSSO_M38_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M39 N_PAD_M40_d N_U28_U42_r1_M39_g N_VSSO_M39_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M40 N_PAD_M40_d N_U28_U42_r1_M40_g N_VSSO_M37_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M35 N_PAD_M41_d N_U15_ngate_M35_g N_VSSO_M35_s N_VSSO_M38_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M41 N_PAD_M41_d N_U28_U42_r1_M41_g N_VSSO_M39_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M31 N_PAD_M36_d N_U17_ngate2_M31_g N_VSSO_M31_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M36 N_PAD_M36_d N_U15_ngate_M36_g N_VSSO_M35_s N_VSSO_M38_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M33 N_PAD_M32_d N_U28_ngate3_M33_g N_VSSO_M33_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M32 N_PAD_M32_d N_U17_ngate2_M32_g N_VSSO_M31_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M42 N_PAD_M34_d N_U28_U42_r1_M42_g N_VSSO_M42_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M34 N_PAD_M34_d N_U28_ngate3_M34_g N_VSSO_M33_s N_VSSO_M38_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M69 N_U28_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M63_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
M56 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56_g N_U28_U72_pgate_M56_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M56@2 N_U15_pgate_M56_d N_net_m56_VSSO_res_M56@2_g N_U28_U72_pgate_M56@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@3 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@3_g N_U28_U72_pgate_M56@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@4 N_U15_pgate_M56@3_d N_net_m56_VSSO_res_M56@4_g N_U28_U72_pgate_M56@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M56@5 N_U15_pgate_M56@5_d N_net_m56_VSSO_res_M56@5_g N_U28_U72_pgate_M56@4_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR61 N_U28_U42_r1_R61_pos N_VSSO_R61_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VSSO_res_RM69_pos N_VSSO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR57 N_noxref_2_R57_pos N_PAD_R57_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR58 N_noxref_2_R58_pos N_U28_padr_R58_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M49 N_VDDO_M49_d N_U28_U71_UN_P_TOP_M49_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M50 N_VDDO_M51_d N_U28_U71_UN_P_TOP_M50_g N_PAD_M49_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M43 N_VDDO_M48_d N_U28_U72_pgate_M43_g N_PAD_M43_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M44 N_VDDO_M44_d N_U28_U72_pgate_M44_g N_PAD_M43_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M51 N_VDDO_M51_d N_U28_U71_UN_P_TOP_M51_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M52 N_VDDO_M52_d N_U28_U71_UN_P_TOP_M52_g N_PAD_M51_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M53 N_VDDO_M52_d N_U28_U71_UN_P_TOP_M53_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M54 N_VDDO_M54_d N_U28_U71_UN_P_TOP_M54_g N_PAD_M53_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M45 N_VDDO_M54_d N_U28_U72_pgate_M45_g N_PAD_M45_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M46 N_VDDO_M46_d N_U28_U72_pgate_M46_g N_PAD_M45_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M47 N_VDDO_M46_d N_U28_U72_pgate_M47_g N_PAD_M47_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M48 N_VDDO_M48_d N_U28_U72_pgate_M48_g N_PAD_M47_s N_VDDO_M51_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M55 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55_g N_U28_U72_pgate_M55_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M55@2 N_U15_pgate_M55_d N_net_m55_VDDO_res_M55@2_g N_U28_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M55@3 N_U15_pgate_M55@3_d N_net_m55_VDDO_res_M55@3_g N_U28_U72_pgate_M55@2_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M62 N_VDDO_M62_d N_net_m62_VDDO_res_M62_g N_U28_U71_UN_P_TOP_M62_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M55_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U15_ngate_M1_g N_VSSO_M1_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M60 N_U28_ngate3_M60_d N_U17_ngatex_M60_g N_VSSO_M60_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U28_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U28_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U30_MPI1_drain_M68_d N_U28_padr_M68_g N_VSSO_M68_s N_VSS_M55_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M28 N_U15_U12_oenb_M28_d N_U15_U15_OUTSHIFT_M28_g N_VSSO_M28_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M7 N_U15_ngate_M7_d N_U15_ISHF_M7_g N_VSSO_M7_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M7@2 N_U15_ngate_M7_d N_U15_ISHF_M7@2_g N_VSSO_M7@2_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M27 N_U15_ngate_M27_d N_U15_U15_OUTSHIFT_M27_g N_VSSO_M7@2_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M8 N_U15_pgate_M8_d N_U15_U12_oenb_M8_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M8@2 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@2_g N_U15_ngate_M8_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M8@3 N_U15_pgate_M8@2_d N_U15_U12_oenb_M8@3_g N_U15_ngate_M8@3_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M21 N_U15_U15_MPLL1_dr_M21_d N_OEN_M21_g N_VSSO_M21_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M23 N_VDDO_M23_d N_U15_U15_MN1_drai_M23_g N_U15_U15_MPLL1_dr_M23_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M21@2 N_U15_U15_MPLL1_dr_M21@2_d N_OEN_M21@2_g N_VSSO_M21_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22 N_U15_U15_OUTSHIFT_M22_d N_U15_U15_MN1_drai_M22_g N_VSSO_M22_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M22@2 N_U15_U15_OUTSHIFT_M22@2_d N_U15_U15_MN1_drai_M22@2_g N_VSSO_M22_s
+ N_VSS_M55_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M15 N_VDDO_M15_d N_U15_U14_MN1_drai_M15_g N_U15_U14_MPLL1_dr_M15_s N_VSS_M55_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M13 N_U15_U14_MPLL1_dr_M13_d N_I_M13_g N_VSSO_M13_s N_VSS_M55_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M13@2 N_U15_U14_MPLL1_dr_M13@2_d N_I_M13@2_g N_VSSO_M13_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14 N_U15_ISHF_M14_d N_U15_U14_MN1_drai_M14_g N_VSSO_M14_s N_VSS_M55_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M14@2 N_U15_ISHF_M14@2_d N_U15_U14_MN1_drai_M14@2_g N_VSSO_M14_s N_VSS_M55_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M16 N_U15_U14_MN1_drai_M16_d N_I_M16_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M24 N_U15_U15_MN1_drai_M24_d N_OEN_M24_g N_VSS_M16_s N_VSS_M55_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M63 N_U28_U71_UN_P_TOP_M63_d N_net_m63_VSSO_res_M63_g N_VDDO_M63_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M63_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M63_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U15_ngate_M2_g N_VDDO_M2_s N_VDDO_M63_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M59 N_U28_ngate3_M59_d N_U17_ngatex_M59_g N_U17_ngate2_M59_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U28_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U30_MPI2_drain N_U28_padr_M64_g N_VDDO_M64_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U30_MPI1_drain_M65_d N_U28_padr_M65_g U30_MPI2_drain N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M29 N_U15_U12_oenb_M29_d N_U15_U15_OUTSHIFT_M29_g N_VDDO_M29_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M29@2 N_U15_U12_oenb_M29@2_d N_U15_U15_OUTSHIFT_M29@2_g N_VDDO_M29_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M9 N_U15_pgate_M9_d N_U15_ISHF_M9_g N_VDDO_M9_s N_VDDO_M63_b PHV L=3.6e-07
+ W=2e-05 AD=1.28e-11 AS=8.2e-12 PD=4.128e-05 PS=2.082e-05
M9@2 N_U15_pgate_M9@2_d N_U15_ISHF_M9@2_g N_VDDO_M9_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=2e-05 AD=9.6e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M30 N_U15_pgate_M9@2_d N_U15_U12_oenb_M30_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=4.8e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M30@2 N_U15_pgate_M30@2_d N_U15_U12_oenb_M30@2_g N_VDDO_M30_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=1e-05 AD=6.3e-12 AS=4.1e-12 PD=2.126e-05 PS=1.082e-05
M10 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10_g N_U15_pgate_M10_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M10@2 N_U15_ngate_M10_d N_U15_U15_OUTSHIFT_M10@2_g N_U15_pgate_M10@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M10@3 N_U15_ngate_M10@3_d N_U15_U15_OUTSHIFT_M10@3_g N_U15_pgate_M10@2_s
+ N_VDDO_M63_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M19 N_U15_U15_MPLL1_dr_M19_d N_U15_U15_OUTSHIFT_M19_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M20 N_U15_U15_OUTSHIFT_M20_d N_U15_U15_MPLL1_dr_M20_g N_VDDO_M19_s N_VDDO_M63_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M11 N_U15_U14_MPLL1_dr_M11_d N_U15_ISHF_M11_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M12 N_U15_ISHF_M12_d N_U15_U14_MPLL1_dr_M12_g N_VDDO_M11_s N_VDDO_M63_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M17 N_U15_U14_MN1_drai_M17_d N_I_M17_g N_VDD_M17_s N_VDD_M17_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M17@2 N_U15_U14_MN1_drai_M17_d N_I_M17@2_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25 N_U15_U15_MN1_drai_M25_d N_OEN_M25_g N_VDD_M17@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M25@2 N_U15_U15_MN1_drai_M25_d N_OEN_M25@2_g N_VDD_M25@2_s N_VDD_M17_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D18 N_VSS_M55_b N_I_D18_neg DN18  AREA=2.5e-13 PJ=2e-06
D26 N_VSS_M55_b N_OEN_D26_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM63 N_VSSO_RM63_pos N_net_m63_VSSO_res_RM63_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM55 N_VDDO_RM55_pos N_net_m55_VDDO_res_RM55_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM62 N_VDDO_RM62_pos N_net_m62_VDDO_res_RM62_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM56 N_net_m56_VSSO_res_RM56_pos N_VSSO_RM56_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359732f
c_2 U30_MPI2_drain 0 0.0169448f
*
.include "pt3t02u.dist.sp.PT3T02U.pxi"
*
.ends
*
*
* File: pt3t03d.dist.sp
* Created: Sun Jul  4 13:11:22 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t03d.dist.sp.pex"
.subckt pt3t03d  PAD I OEN VDD VSS VDDO VSSO 
* 
M69 N_U29_padr_M69_d N_net_m69_VDDO_res_M69_g U31_U22_source N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=1.56e-12 AS=4e-13 PD=5.56e-06 PS=2.4e-06
M70 U31_U22_source N_net_m70_VDDO_res_M70_g N_VSSO_M70_s N_VSS_M19_b NHV
+ L=5.5e-06 W=2e-06 AD=4e-13 AS=1.56e-12 PD=2.4e-06 PS=5.56e-06
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_net_m69_VDDO_res_RM69_pos N_VDDO_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM70 N_VDDO_RM69_neg N_net_m70_VDDO_res_RM70_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U32_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U32_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U32_MPI1_drain_M65_d N_U29_padr_M65_g U32_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U32_MPI2_drain 0 0.0169448f
*
.include "pt3t03d.dist.sp.PT3T03D.pxi"
*
.ends
*
*
* File: pt3t03.dist.sp
* Created: Sun Jul  4 13:09:47 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t03.dist.sp.pex"
.subckt pt3t03  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U31_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U31_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U31_MPI1_drain_M65_d N_U29_padr_M65_g U31_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U31_MPI2_drain 0 0.0169448f
*
.include "pt3t03.dist.sp.PT3T03.pxi"
*
.ends
*
*
* File: pt3t03u.dist.sp
* Created: Sun Jul  4 13:11:28 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pt3t03u.dist.sp.pex"
.subckt pt3t03u  PAD I OEN VDD VSS VDDO VSSO 
* 
M15 N_PAD_M13_d N_U30_ngate_M15_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M13 N_PAD_M13_d N_U29_U42_r1_M13_g N_VSSO_M13_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M16 N_PAD_M17_d N_U30_ngate_M16_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M17 N_PAD_M17_d N_U30_ngate_M17_g N_VSSO_M15_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M9 N_PAD_M18_d N_U17_ngate2_M9_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M18 N_PAD_M18_d N_U30_ngate_M18_g N_VSSO_M16_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M10 N_PAD_M11_d N_U17_ngate2_M10_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M11 N_PAD_M11_d N_U17_ngate2_M11_g N_VSSO_M9_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M7 N_PAD_M12_d N_U29_ngate3_M7_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M12 N_PAD_M12_d N_U17_ngate2_M12_g N_VSSO_M10_s N_VSSO_M13_b NHV L=5e-07
+ W=3e-05 AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M14 N_PAD_M8_d N_U29_U42_r1_M14_g N_VSSO_M14_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=3.99e-11 PD=3.672e-05 PS=6.266e-05
M8 N_PAD_M8_d N_U29_ngate3_M8_g N_VSSO_M7_s N_VSSO_M13_b NHV L=5e-07 W=3e-05
+ AD=1.008e-10 AS=2.58e-11 PD=3.672e-05 PS=3.172e-05
M20 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20_g N_U29_U72_pgate_M20_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M20@2 N_U30_pgate_M20_d N_net_m20_VSSO_res_M20@2_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@3 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@3_g N_U29_U72_pgate_M20@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@4 N_U30_pgate_M20@3_d N_net_m20_VSSO_res_M20@4_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M20@5 N_U30_pgate_M20@5_d N_net_m20_VSSO_res_M20@5_g N_U29_U72_pgate_M20@4_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M69 N_U29_padr_M69_d N_net_m69_VSSO_res_M69_g N_VDDO_M69_s N_VDDO_M39_b PHV
+ L=2e-06 W=2e-06 AD=4e-12 AS=4e-12 PD=8e-06 PS=8e-06
XR37 N_U29_U42_r1_R37_pos N_VSSO_R37_neg RNWELLSTI2T w=2.1e-06 l=8.65e-06 
XRM69 N_VSSO_RM69_pos N_net_m69_VSSO_res_RM69_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XR21 N_noxref_2_R21_pos N_PAD_R21_neg RNMPOLY2T w=4e-06 l=2.5e-06 
XR22 N_noxref_2_R22_pos N_U29_padr_R22_neg RNMPOLY2T w=4e-06 l=2.5e-06 
M35 N_VDDO_M35_d N_U29_U71_UN_P_TOP_M35_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M36 N_VDDO_M27_d N_U29_U71_UN_P_TOP_M36_g N_PAD_M35_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M25 N_VDDO_M34_d N_U29_U72_pgate_M25_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M26 N_VDDO_M26_d N_U29_U72_pgate_M26_g N_PAD_M25_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=7.384e-11 AS=1.2064e-10 PD=0.00010684 PS=5.664e-05
M27 N_VDDO_M27_d N_U29_U72_pgate_M27_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M28 N_VDDO_M28_d N_U29_U72_pgate_M28_g N_PAD_M27_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M29 N_VDDO_M28_d N_U29_U72_pgate_M29_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M30 N_VDDO_M30_d N_U29_U72_pgate_M30_g N_PAD_M29_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M31 N_VDDO_M30_d N_U29_U72_pgate_M31_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M32 N_VDDO_M32_d N_U29_U72_pgate_M32_g N_PAD_M31_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M33 N_VDDO_M32_d N_U29_U72_pgate_M33_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M34 N_VDDO_M34_d N_U29_U72_pgate_M34_g N_PAD_M33_s N_VDDO_M27_b PHV L=4e-07
+ W=5.2e-05 AD=4.732e-11 AS=1.2064e-10 PD=5.382e-05 PS=5.664e-05
M19 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19_g N_U29_U72_pgate_M19_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=1.03354e-11 PD=1.749e-05
+ PS=3.458e-05
M19@2 N_U30_pgate_M19_d N_net_m19_VDDO_res_M19@2_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=6.8347e-12 AS=6.8347e-12 PD=1.749e-05
+ PS=1.749e-05
M19@3 N_U30_pgate_M19@3_d N_net_m19_VDDO_res_M19@3_g N_U29_U72_pgate_M19@2_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1.667e-05 AD=1.05021e-11 AS=6.8347e-12 PD=3.46e-05
+ PS=1.749e-05
M38 N_VDDO_M38_d N_net_m38_VDDO_res_M38_g N_U29_U71_UN_P_TOP_M38_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M3 N_U17_ngate2_M3_d N_I_M3_g N_VSSO_M3_s N_VSS_M19_b NHV L=3.6e-07 W=1.5e-05
+ AD=9.3e-12 AS=9.3e-12 PD=3.124e-05 PS=3.124e-05
M4 N_U17_ngate2_M4_d N_U17_ngatex_M4_g N_VSSO_M4_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-06 AD=6.2e-13 AS=6.2e-13 PD=3.24e-06 PS=3.24e-06
M1 N_U17_ngatex_M1_d N_U30_ngate_M1_g N_VSSO_M1_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M24 N_U29_ngate3_M24_d N_U17_ngatex_M24_g N_VSSO_M24_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M67 N_U29_padr_M67_d N_net_m67_VSSO_res_M67_g N_VSSO_M67_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M67@2 N_U29_padr_M67@2_d N_net_m67_VSSO_res_M67@2_g N_VSSO_M67_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M68 N_U32_MPI1_drain_M68_d N_U29_padr_M68_g N_VSSO_M68_s N_VSS_M19_b NHV
+ L=3.6e-07 W=6e-06 AD=3.72e-12 AS=3.72e-12 PD=1.324e-05 PS=1.324e-05
M61 N_U30_U12_oenb_M61_d N_U30_U15_OUTSHIFT_M61_g N_VSSO_M61_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=6.2e-12 PD=2.124e-05 PS=2.124e-05
M42 N_U30_ngate_M42_d N_U30_ISHF_M42_g N_VSSO_M42_s N_VSS_M19_b NHV L=3.6e-07
+ W=1.5e-05 AD=6.15e-12 AS=9.3e-12 PD=1.582e-05 PS=3.124e-05
M42@2 N_U30_ngate_M42_d N_U30_ISHF_M42@2_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.5e-05 AD=6.15e-12 AS=6.97793e-12 PD=1.582e-05 PS=1.89385e-05
M60 N_U30_ngate_M60_d N_U30_U15_OUTSHIFT_M60_g N_VSSO_M42@2_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1.006e-05 AD=6.2372e-12 AS=4.67987e-12 PD=2.136e-05 PS=1.27015e-05
M43 N_U30_pgate_M43_d N_U30_U12_oenb_M43_g N_U30_ngate_M43_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M43@2 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@2_g N_U30_ngate_M43_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05 PS=1.082e-05
M43@3 N_U30_pgate_M43@2_d N_U30_U12_oenb_M43@3_g N_U30_ngate_M43@3_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05
+ PS=2.124e-05
M54 N_U30_U15_MPLL1_dr_M54_d N_OEN_M54_g N_VSSO_M54_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.6e-12 AS=4.1e-12 PD=2.132e-05 PS=1.082e-05
M56 N_VDDO_M56_d N_U30_U15_MN1_drai_M56_g N_U30_U15_MPLL1_dr_M56_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M54@2 N_U30_U15_MPLL1_dr_M54@2_d N_OEN_M54@2_g N_VSSO_M54_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55 N_U30_U15_OUTSHIFT_M55_d N_U30_U15_MN1_drai_M55_g N_VSSO_M55_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M55@2 N_U30_U15_OUTSHIFT_M55@2_d N_U30_U15_MN1_drai_M55@2_g N_VSSO_M55_s
+ N_VSS_M19_b NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M48 N_VDDO_M48_d N_U30_U14_MN1_drai_M48_g N_U30_U14_MPLL1_dr_M48_s N_VSS_M19_b
+ NHV L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M46 N_U30_U14_MPLL1_dr_M46_d N_I_M46_g N_VSSO_M46_s N_VSS_M19_b NHV L=3.6e-07
+ W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M46@2 N_U30_U14_MPLL1_dr_M46@2_d N_I_M46@2_g N_VSSO_M46_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47 N_U30_ISHF_M47_d N_U30_U14_MN1_drai_M47_g N_VSSO_M47_s N_VSS_M19_b NHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M47@2 N_U30_ISHF_M47@2_d N_U30_U14_MN1_drai_M47@2_g N_VSSO_M47_s N_VSS_M19_b
+ NHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M49 N_U30_U14_MN1_drai_M49_d N_I_M49_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.925e-12 AS=1.8375e-12 PD=1.117e-05 PS=5.735e-06
M57 N_U30_U15_MN1_drai_M57_d N_OEN_M57_g N_VSS_M49_s N_VSS_M19_b N18 L=1.8e-07
+ W=5e-06 AD=2.9e-12 AS=1.8375e-12 PD=1.116e-05 PS=5.735e-06
M39 N_U29_U71_UN_P_TOP_M39_d N_net_m39_VSSO_res_M39_g N_VDDO_M39_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M6 U17_U15_U8_sourc N_I_M6_g N_VDDO_M6_s N_VDDO_M39_b PHV L=3.6e-07 W=1.5e-05
+ AD=3.45e-12 AS=9.3e-12 PD=1.546e-05 PS=3.124e-05
M5 N_U17_ngate2_M5_d N_U17_ngatex_M5_g U17_U15_U8_sourc N_VDDO_M39_b PHV
+ L=3.6e-07 W=1.5e-05 AD=1.02e-11 AS=3.45e-12 PD=3.136e-05 PS=1.546e-05
M2 N_U17_ngatex_M2_d N_U30_ngate_M2_g N_VDDO_M2_s N_VDDO_M39_b PHV L=3.6e-07
+ W=7e-06 AD=4.34e-12 AS=4.34e-12 PD=1.524e-05 PS=1.524e-05
M23 N_U29_ngate3_M23_d N_U17_ngatex_M23_g N_U17_ngate2_M23_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=5e-06 AD=3.1e-12 AS=3.1e-12 PD=1.124e-05 PS=1.124e-05
M66 N_U29_padr_M66_d N_net_m66_VDDO_res_M66_g N_VDDO_M66_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=1.24e-11 PD=4.124e-05 PS=4.124e-05
M64 U32_MPI2_drain N_U29_padr_M64_g N_VDDO_M64_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=4e-12 AS=1.24e-11 PD=2.04e-05 PS=4.124e-05
M65 N_U32_MPI1_drain_M65_d N_U29_padr_M65_g U32_MPI2_drain N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=1.24e-11 AS=4e-12 PD=4.124e-05 PS=2.04e-05
M62 N_U30_U12_oenb_M62_d N_U30_U15_OUTSHIFT_M62_g N_VDDO_M62_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M62@2 N_U30_U12_oenb_M62@2_d N_U30_U15_OUTSHIFT_M62@2_g N_VDDO_M62_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05
+ PS=1.082e-05
M40 N_U30_pgate_M40_d N_U30_ISHF_M40_g N_VDDO_M40_s N_VDDO_M39_b PHV L=3.6e-07
+ W=2e-05 AD=8.2e-12 AS=1.24e-11 PD=2.082e-05 PS=4.124e-05
M40@2 N_U30_pgate_M40_d N_U30_ISHF_M40@2_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=8.2e-12 AS=8.2e-12 PD=2.082e-05 PS=2.082e-05
M40@3 N_U30_pgate_M40@3_d N_U30_ISHF_M40@3_g N_VDDO_M40@2_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=2e-05 AD=9.66667e-12 AS=8.2e-12 PD=2.776e-05 PS=2.082e-05
M63 N_U30_pgate_M40@3_d N_U30_U12_oenb_M63_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=4.83333e-12 AS=4.1e-12 PD=1.388e-05 PS=1.082e-05
M63@2 N_U30_pgate_M63@2_d N_U30_U12_oenb_M63@2_g N_VDDO_M63_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=1e-05 AD=6.2e-12 AS=4.1e-12 PD=2.124e-05 PS=1.082e-05
M41 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41_g N_U30_pgate_M41_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=6.2e-12 PD=1.082e-05 PS=2.124e-05
M41@2 N_U30_ngate_M41_d N_U30_U15_OUTSHIFT_M41@2_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=4.1e-12 AS=4.1e-12 PD=1.082e-05
+ PS=1.082e-05
M41@3 N_U30_ngate_M41@3_d N_U30_U15_OUTSHIFT_M41@3_g N_U30_pgate_M41@2_s
+ N_VDDO_M39_b PHV L=3.6e-07 W=1e-05 AD=7.2e-12 AS=4.1e-12 PD=2.144e-05
+ PS=1.082e-05
M52 N_U30_U15_MPLL1_dr_M52_d N_U30_U15_OUTSHIFT_M52_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M53 N_U30_U15_OUTSHIFT_M53_d N_U30_U15_MPLL1_dr_M53_g N_VDDO_M52_s N_VDDO_M39_b
+ PHV L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M44 N_U30_U14_MPLL1_dr_M44_d N_U30_ISHF_M44_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M45 N_U30_ISHF_M45_d N_U30_U14_MPLL1_dr_M45_g N_VDDO_M44_s N_VDDO_M39_b PHV
+ L=3.6e-07 W=7.2e-06 AD=4.464e-12 AS=2.952e-12 PD=1.564e-05 PS=8.02e-06
M50 N_U30_U14_MN1_drai_M50_d N_I_M50_g N_VDD_M50_s N_VDD_M50_b P18 L=1.8e-07
+ W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
M50@2 N_U30_U14_MN1_drai_M50_d N_I_M50@2_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58 N_U30_U15_MN1_drai_M58_d N_OEN_M58_g N_VDD_M50@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=1.4e-12 PD=5.56e-06 PS=5.56e-06
M58@2 N_U30_U15_MN1_drai_M58_d N_OEN_M58@2_g N_VDD_M58@2_s N_VDD_M50_b P18
+ L=1.8e-07 W=5e-06 AD=1.4e-12 AS=2.45e-12 PD=5.56e-06 PS=1.098e-05
D51 N_VSS_M19_b N_I_D51_neg DN18  AREA=2.5e-13 PJ=2e-06
D59 N_VSS_M19_b N_OEN_D59_neg DN18  AREA=2.5e-13 PJ=2e-06
XRM39 N_VSSO_RM39_pos N_net_m39_VSSO_res_RM39_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM66 N_net_m66_VDDO_res_RM66_pos N_VDDO_RM66_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM19 N_VDDO_RM19_pos N_net_m19_VDDO_res_RM19_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM38 N_VDDO_RM38_pos N_net_m38_VDDO_res_RM38_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM67 N_VSSO_RM67_pos N_net_m67_VSSO_res_RM67_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
XRM20 N_net_m20_VSSO_res_RM20_pos N_VSSO_RM20_neg RPMPOLY2T w=2e-06 l=6.455e-06
+ 
c_1 U17_U15_U8_sourc 0 0.359751f
c_2 U32_MPI2_drain 0 0.0169448f
*
.include "pt3t03u.dist.sp.PT3T03U.pxi"
*
.ends
*
*
* File: pv0a.dist.sp
* Created: Sun Jul  4 13:13:09 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0a.dist.sp.pex"
.subckt pv0a  VSSO VDD VSS VDDO 
* 
M4 N_VDDO_M5_d N_U31_U29_c2_M4_g N_VSSO_M11_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDO_M5_d N_U31_U29_c2_M5_g N_VSSO_M5_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDO_M7_d N_U31_U29_c2_M6_g N_VSSO_M6_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M7 N_VDDO_M7_d N_U31_U29_c2_M7_g N_VSSO_M12_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDO_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U19_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U31_U29_c2_R2_pos N_noxref_6_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_6_R3_pos N_VSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M8 N_VDDO_M8_d N_U31_U29_c2_M8_g N_VSSO_M8_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M9 N_VDDO_M8_d N_U31_U29_c2_M9_g N_VSSO_M9_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M10 N_VDDO_M10_d N_U31_U29_c2_M10_g N_VSSO_M9_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDO_M10_d N_U31_U29_c2_M11_g N_VSSO_M11_s N_VSSO_M8_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDO_M12_d N_U31_U29_c2_M12_g N_VSSO_M12_s N_VSSO_M8_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDO_M12_d N_U31_U29_c2_M13_g N_VSSO_M13_s N_VSSO_M8_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDO_M14_d N_U31_U29_c2_M14_g N_VSSO_M13_s N_VSSO_M8_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDO_M14_d N_U31_U29_c2_M15_g N_VSSO_M8_s N_VSSO_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
D31@2 N_VSSO_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSSO_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSSO_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSSO_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSSO_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSSO_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSSO_D31@8_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSSO_D31@9_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSSO_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@2 N_VSS_D30@2_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSS_D30@3_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSS_D30@4_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSS_D30@5_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSS_D30@6_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSS_D30@7_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSS_D30@8_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSS_D30@9_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSS_D30_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC4_5 N_VDDO_C4_5_pos N_U31_U29_c2_C4_5_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSSO_M16_d N_U19_U22$11_gate_M16_g N_VDDO_M16_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSSO_M16_d N_U19_U22$11_gate_M17_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSSO_M18_d N_U19_U22$11_gate_M18_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSSO_M18_d N_U19_U22$11_gate_M19_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSSO_M20_d N_U19_U22$11_gate_M20_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSSO_M20_d N_U19_U22$11_gate_M21_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSSO_M22_d N_U19_U22$11_gate_M22_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSSO_M22_d N_U19_U22$11_gate_M23_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSSO_M24_d N_U19_U22$11_gate_M24_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSSO_M24_d N_U19_U22$11_gate_M25_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSSO_M26_d N_U19_U22$11_gate_M26_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSSO_M26_d N_U19_U22$11_gate_M27_g N_VDDO_M27_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pv0a.dist.sp.PV0A.pxi"
*
.ends
*
*
* File: pv0c.dist.sp
* Created: Sun Jul  4 13:13:03 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0c.dist.sp.pex"
.subckt pv0c  VSSC VDD VSS VDDO VSSO 
* 
M18 N_VDD_M19_d N_U33_U29_c2_M18_g N_VSSC_M25_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_VDD_M19_d N_U33_U29_c2_M19_g N_VSSC_M19_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_VDD_M21_d N_U33_U29_c2_M20_g N_VSSC_M20_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M21 N_VDD_M21_d N_U33_U29_c2_M21_g N_VSSC_M26_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_VDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U34_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_U33_U29_c2_R16_pos N_noxref_7_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR17 N_noxref_7_R17_pos N_VSSC_R17_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M22 N_VDD_M22_d N_U33_U29_c2_M22_g N_VSSC_M22_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M23 N_VDD_M22_d N_U33_U29_c2_M23_g N_VSSC_M23_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M24 N_VDD_M24_d N_U33_U29_c2_M24_g N_VSSC_M23_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_VDD_M24_d N_U33_U29_c2_M25_g N_VSSC_M25_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_VDD_M26_d N_U33_U29_c2_M26_g N_VSSC_M26_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_VDD_M26_d N_U33_U29_c2_M27_g N_VSSC_M27_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_VDD_M28_d N_U33_U29_c2_M28_g N_VSSC_M27_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_VDD_M28_d N_U33_U29_c2_M29_g N_VSSC_M22_s N_VSSC_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M3 N_VSSC_M3_d N_U34_U31_r2_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
M4 N_VSSC_M3_d N_U34_U31_r2_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M5 N_VSSC_M5_d N_U34_U31_r2_M5_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M6 N_VSSC_M5_d N_U34_U31_r2_M6_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M7 N_VSSC_M7_d N_U34_U31_r2_M7_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M8 N_VSSC_M7_d N_U34_U31_r2_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M9 N_VSSC_M9_d N_U34_U31_r2_M9_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M10 N_VSSC_M9_d N_U34_U31_r2_M10_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M11 N_VSSC_M11_d N_U34_U31_r2_M11_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M12 N_VSSC_M11_d N_U34_U31_r2_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M13 N_VSSC_M13_d N_U34_U31_r2_M13_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M14 N_VSSC_M13_d N_U34_U31_r2_M14_g N_VDD_M14_s N_VDD_M3_b P18 L=2.5e-07
+ W=4e-05 AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
D30@2 N_VSSC_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSSC_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSSC_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSSC_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSSC_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSSC_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSSC_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSSC_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSSC_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_VSSC_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC8_1 N_VDD_C8_1_pos N_U33_U29_c2_C8_1_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "pv0c.dist.sp.PV0C.pxi"
*
.ends
*
*
* File: pv0f.dist.sp
* Created: Sun Jul  4 13:14:38 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0f.dist.sp.pex"
.subckt pv0f  VSS VDD VDDO VSSO 
* 
M4 N_VDDO_M5_d N_U37_U29_c2_M4_g N_VSS_M11_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDO_M5_d N_U37_U29_c2_M5_g N_VSS_M5_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDO_M7_d N_U37_U29_c2_M6_g N_VSS_M6_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M7 N_VDDO_M7_d N_U37_U29_c2_M7_g N_VSS_M12_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDO_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U34_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U37_U29_c2_R2_pos N_noxref_6_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_6_R3_pos N_VSS_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M8 N_VDDO_M8_d N_U37_U29_c2_M8_g N_VSS_M8_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M9 N_VDDO_M8_d N_U37_U29_c2_M9_g N_VSS_M9_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M10 N_VDDO_M10_d N_U37_U29_c2_M10_g N_VSS_M9_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDO_M10_d N_U37_U29_c2_M11_g N_VSS_M11_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDO_M12_d N_U37_U29_c2_M12_g N_VSS_M12_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDO_M12_d N_U37_U29_c2_M13_g N_VSS_M13_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDO_M14_d N_U37_U29_c2_M14_g N_VSS_M13_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDO_M14_d N_U37_U29_c2_M15_g N_VSS_M8_s N_VSS_M8_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
dX23/D0_noxref N_VSS_X23/D0_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D1_noxref N_VSS_X23/D1_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D2_noxref N_VSS_X23/D2_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D3_noxref N_VSS_X23/D3_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D4_noxref N_VSS_X23/D4_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D5_noxref N_VSS_X23/D5_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D6_noxref N_VSS_X23/D6_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D7_noxref N_VSS_X23/D7_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D8_noxref N_VSS_X23/D8_noxref_pos N_VSS_X23/D0_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D9_noxref N_VSS_X23/D9_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D10_noxref N_VSS_X23/D10_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D11_noxref N_VSS_X23/D11_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D12_noxref N_VSS_X23/D12_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D13_noxref N_VSS_X23/D13_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D14_noxref N_VSS_X23/D14_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D15_noxref N_VSS_X23/D15_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D16_noxref N_VSS_X23/D16_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
dX23/D17_noxref N_VSS_X23/D17_noxref_pos N_VSS_X23/D9_noxref_neg DPH 
+ AREA=1.331e-11 PJ=2.862e-05
XC3_5 N_VDDO_C3_5_pos N_U37_U29_c2_C3_5_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSS_M16_d N_U34_U22$11_gate_M16_g N_VDDO_M16_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSS_M16_d N_U34_U22$11_gate_M17_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSS_M18_d N_U34_U22$11_gate_M18_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSS_M18_d N_U34_U22$11_gate_M19_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSS_M20_d N_U34_U22$11_gate_M20_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSS_M20_d N_U34_U22$11_gate_M21_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSS_M22_d N_U34_U22$11_gate_M22_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSS_M22_d N_U34_U22$11_gate_M23_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSS_M24_d N_U34_U22$11_gate_M24_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSS_M24_d N_U34_U22$11_gate_M25_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSS_M26_d N_U34_U22$11_gate_M26_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSS_M26_d N_U34_U22$11_gate_M27_g N_VDDO_M27_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pv0f.dist.sp.PV0F.pxi"
*
.ends
*
*
* File: pv0i.dist.sp
* Created: Sun Jul  4 13:14:33 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pv0i.dist.sp.pex"
.subckt pv0i  VSS VDD VDDO VSSO 
* 
M18 N_VDD_M19_d N_U31_U18_r1_M18_g N_VSS_M25_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_VDD_M19_d N_U31_U18_r1_M19_g N_VSS_M19_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_VDD_M21_d N_U31_U18_r1_M20_g N_VSS_M20_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M21 N_VDD_M21_d N_U31_U18_r1_M21_g N_VSS_M26_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_VDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U33_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR15 N_U31_U18_r1_R15_pos N_noxref_6_R15_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_noxref_6_R16_pos N_VSS_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M22 N_VDD_M22_d N_U31_U18_r1_M22_g N_VSS_M22_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M23 N_VDD_M22_d N_U31_U18_r1_M23_g N_VSS_M23_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M24 N_VDD_M24_d N_U31_U18_r1_M24_g N_VSS_M23_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_VDD_M24_d N_U31_U18_r1_M25_g N_VSS_M25_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_VDD_M26_d N_U31_U18_r1_M26_g N_VSS_M26_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_VDD_M26_d N_U31_U18_r1_M27_g N_VSS_M27_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_VDD_M28_d N_U31_U18_r1_M28_g N_VSS_M27_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_VDD_M28_d N_U31_U18_r1_M29_g N_VSS_M22_s N_VSS_M22_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M3 N_VSS_M3_d N_U33_U31_r2_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
M4 N_VSS_M3_d N_U33_U31_r2_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M5 N_VSS_M5_d N_U33_U31_r2_M5_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M6 N_VSS_M5_d N_U33_U31_r2_M6_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M7 N_VSS_M7_d N_U33_U31_r2_M7_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M8 N_VSS_M7_d N_U33_U31_r2_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M9 N_VSS_M9_d N_U33_U31_r2_M9_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M10 N_VSS_M9_d N_U33_U31_r2_M10_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M11 N_VSS_M11_d N_U33_U31_r2_M11_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M12 N_VSS_M11_d N_U33_U31_r2_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M13 N_VSS_M13_d N_U33_U31_r2_M13_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M14 N_VSS_M13_d N_U33_U31_r2_M14_g N_VDD_M14_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
D30@2 N_VSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC8_1 N_VDD_C8_1_pos N_U31_U18_r1_C8_1_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "pv0i.dist.sp.PV0I.pxi"
*
.ends
*
*
* File: pvda.dist.sp
* Created: Sun Jul  4 13:18:02 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pvda.dist.sp.pex"
.subckt pvda  VDDO VDD VSS VSSO 
* 
M4 N_VDDO_M10_d N_U30_U29_c2_M4_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDO_M11_d N_U30_U29_c2_M5_g N_VSSO_M5_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDO_M12_d N_U30_U29_c2_M6_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_VDDO_M13_d N_U30_U29_c2_M7_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_VDDO_M14_d N_U30_U29_c2_M8_g N_VSSO_M8_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_VDDO_M15_d N_U30_U29_c2_M9_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDO_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U19_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U30_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_VSSO_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_VDDO_M10_d N_U30_U29_c2_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDO_M11_d N_U30_U29_c2_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDO_M12_d N_U30_U29_c2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDO_M13_d N_U30_U29_c2_M13_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDO_M14_d N_U30_U29_c2_M14_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDO_M15_d N_U30_U29_c2_M15_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
D31@2 N_VSSO_D31@2_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSSO_D31@3_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSSO_D31@4_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSSO_D31@5_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSSO_D31@6_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSSO_D31@7_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSSO_D31@8_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSSO_D31@9_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSSO_D31_pos N_VSS_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@2 N_VSS_D30@2_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSS_D30@3_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSS_D30@4_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSS_D30@5_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSS_D30@6_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSS_D30@7_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSS_D30@8_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSS_D30@9_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSS_D30_pos N_VSSO_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC3_5 N_VDDO_C3_5_pos N_U30_U29_c2_C3_5_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSSO_M16_d N_U19_U22$11_gate_M16_g N_VDDO_M16_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSSO_M16_d N_U19_U22$11_gate_M17_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSSO_M18_d N_U19_U22$11_gate_M18_g N_VDDO_M17_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSSO_M18_d N_U19_U22$11_gate_M19_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSSO_M20_d N_U19_U22$11_gate_M20_g N_VDDO_M19_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSSO_M20_d N_U19_U22$11_gate_M21_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSSO_M22_d N_U19_U22$11_gate_M22_g N_VDDO_M21_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSSO_M22_d N_U19_U22$11_gate_M23_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSSO_M24_d N_U19_U22$11_gate_M24_g N_VDDO_M23_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSSO_M24_d N_U19_U22$11_gate_M25_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSSO_M26_d N_U19_U22$11_gate_M26_g N_VDDO_M25_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSSO_M26_d N_U19_U22$11_gate_M27_g N_VDDO_M27_s N_VDDO_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pvda.dist.sp.PVDA.pxi"
*
.ends
*
*
* File: pvdc.dist.sp
* Created: Sun Jul  4 13:17:59 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pvdc.dist.sp.pex"
.subckt pvdc  VDDC VDD VSS VDDO VSSO 
* 
M4 N_VDDC_M10_d N_U36_U29_c2_M4_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M5 N_VDDC_M11_d N_U36_U29_c2_M5_g N_VSSO_M5_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M6 N_VDDC_M12_d N_U36_U29_c2_M6_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M7 N_VDDC_M13_d N_U36_U29_c2_M7_g N_VSSO_M4_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M8 N_VDDC_M14_d N_U36_U29_c2_M8_g N_VSSO_M8_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=3.99e-11 PD=3.692e-05 PS=6.266e-05
M9 N_VDDC_M15_d N_U36_U29_c2_M9_g N_VSSO_M6_s N_VSSO_M10_b NHV L=4e-07 W=3e-05
+ AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
XR28 N_VDDC_R28_pos N_noxref_3_R28_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR29 N_noxref_3_R29_pos N_U35_U22$11_gate_R29_neg RNWELLSTI2T w=2.1e-06
+ l=1.46e-05 
XR2 N_U36_U29_c2_R2_pos N_noxref_5_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR3 N_noxref_5_R3_pos N_VSS_R3_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M10 N_VDDC_M10_d N_U36_U29_c2_M10_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M11 N_VDDC_M11_d N_U36_U29_c2_M11_g N_VSSO_M10_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M12 N_VDDC_M12_d N_U36_U29_c2_M12_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M13 N_VDDC_M13_d N_U36_U29_c2_M13_g N_VSSO_M12_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M14 N_VDDC_M14_d N_U36_U29_c2_M14_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
M15 N_VDDC_M15_d N_U36_U29_c2_M15_g N_VSSO_M14_s N_VSSO_M10_b NHV L=4e-07
+ W=3e-05 AD=1.038e-10 AS=2.58e-11 PD=3.692e-05 PS=3.172e-05
D30@2 N_VSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC3_6 N_VDDC_C3_6_pos N_U36_U29_c2_C3_6_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
M16 N_VSS_M16_d N_U35_U22$11_gate_M16_g N_VDDC_M16_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
M17 N_VSS_M16_d N_U35_U22$11_gate_M17_g N_VDDC_M17_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M18 N_VSS_M18_d N_U35_U22$11_gate_M18_g N_VDDC_M17_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M19 N_VSS_M18_d N_U35_U22$11_gate_M19_g N_VDDC_M19_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M20 N_VSS_M20_d N_U35_U22$11_gate_M20_g N_VDDC_M19_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M21 N_VSS_M20_d N_U35_U22$11_gate_M21_g N_VDDC_M21_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M22 N_VSS_M22_d N_U35_U22$11_gate_M22_g N_VDDC_M21_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M23 N_VSS_M22_d N_U35_U22$11_gate_M23_g N_VDDC_M23_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M24 N_VSS_M24_d N_U35_U22$11_gate_M24_g N_VDDC_M23_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M25 N_VSS_M24_d N_U35_U22$11_gate_M25_g N_VDDC_M25_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M26 N_VSS_M26_d N_U35_U22$11_gate_M26_g N_VDDC_M25_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=3.64e-11 PD=4.464e-05 PS=4.182e-05
M27 N_VSS_M26_d N_U35_U22$11_gate_M27_g N_VDDC_M27_s N_VDDC_M16_b PHV L=4e-07
+ W=4e-05 AD=9.28e-11 AS=5.68e-11 PD=4.464e-05 PS=8.284e-05
*
.include "pvdc.dist.sp.PVDC.pxi"
*
.ends
*
*
* File: pvdi.dist.sp
* Created: Sun Jul  4 13:19:19 2010
* Program "Calibre xRC"
* Version "v2008.4_19.14"
* 
.include "pvdi.dist.sp.pex"
.subckt pvdi  VDD VSS VDDO VSSO 
* 
M18 N_VDD_M24_d N_U31_U18_r1_M18_g N_VSSO_M18_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M19 N_VDD_M25_d N_U31_U18_r1_M19_g N_VSSO_M19_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M20 N_VDD_M26_d N_U31_U18_r1_M20_g N_VSSO_M20_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M21 N_VDD_M27_d N_U31_U18_r1_M21_g N_VSSO_M18_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M22 N_VDD_M28_d N_U31_U18_r1_M22_g N_VSSO_M22_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=3.99e-11 PD=3.722e-05 PS=6.266e-05
M23 N_VDD_M29_d N_U31_U18_r1_M23_g N_VSSO_M20_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
XR1 N_VDD_R1_pos N_noxref_3_R1_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR2 N_noxref_3_R2_pos N_U32_U31_r2_R2_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR15 N_U31_U18_r1_R15_pos N_noxref_5_R15_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
XR16 N_noxref_5_R16_pos N_VSS_R16_neg RNWELLSTI2T w=2.1e-06 l=1.46e-05 
M24 N_VDD_M24_d N_U31_U18_r1_M24_g N_VSSO_M24_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M25 N_VDD_M25_d N_U31_U18_r1_M25_g N_VSSO_M24_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M26 N_VDD_M26_d N_U31_U18_r1_M26_g N_VSSO_M26_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M27 N_VDD_M27_d N_U31_U18_r1_M27_g N_VSSO_M26_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M28 N_VDD_M28_d N_U31_U18_r1_M28_g N_VSSO_M28_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M29 N_VDD_M29_d N_U31_U18_r1_M29_g N_VSSO_M28_s N_VSSO_M24_b N18 L=2.5e-07
+ W=3e-05 AD=1.083e-10 AS=2.58e-11 PD=3.722e-05 PS=3.172e-05
M3 N_VSS_M3_d N_U32_U31_r2_M3_g N_VDD_M3_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
M4 N_VSS_M3_d N_U32_U31_r2_M4_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M5 N_VSS_M5_d N_U32_U31_r2_M5_g N_VDD_M4_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M6 N_VSS_M5_d N_U32_U31_r2_M6_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M7 N_VSS_M7_d N_U32_U31_r2_M7_g N_VDD_M6_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M8 N_VSS_M7_d N_U32_U31_r2_M8_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M9 N_VSS_M9_d N_U32_U31_r2_M9_g N_VDD_M8_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M10 N_VSS_M9_d N_U32_U31_r2_M10_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M11 N_VSS_M11_d N_U32_U31_r2_M11_g N_VDD_M10_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M12 N_VSS_M11_d N_U32_U31_r2_M12_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M13 N_VSS_M13_d N_U32_U31_r2_M13_g N_VDD_M12_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=3.44e-11 PD=4.504e-05 PS=4.172e-05
M14 N_VSS_M13_d N_U32_U31_r2_M14_g N_VDD_M14_s N_VDD_M3_b P18 L=2.5e-07 W=4e-05
+ AD=1.008e-10 AS=5.48e-11 PD=4.504e-05 PS=8.274e-05
D30@2 N_VSSO_D30@2_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@3 N_VSSO_D30@3_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@4 N_VSSO_D30@4_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@5 N_VSSO_D30@5_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@6 N_VSSO_D30@6_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@7 N_VSSO_D30@7_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@8 N_VSSO_D30@8_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30@9 N_VSSO_D30@9_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D30 N_VSSO_D30_pos N_VSS_D30@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@2 N_VSS_D31@2_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@3 N_VSS_D31@3_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@4 N_VSS_D31@4_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@5 N_VSS_D31@5_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@6 N_VSS_D31@6_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@7 N_VSS_D31@7_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@8 N_VSS_D31@8_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31@9 N_VSS_D31@9_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
D31 N_VSS_D31_pos N_VSSO_D31@2_neg DPH  AREA=1.331e-11 PJ=2.862e-05
XC8_1 N_VDD_C8_1_pos N_U31_U18_r1_C8_1_neg NWCAPH2T  L=1.513e-05 W=1.513e-05
*
.include "pvdi.dist.sp.PVDI.pxi"
*
.ends
*
*
